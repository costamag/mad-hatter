module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 ;
  wire n9 , n10 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n22 , n23 , n25 , n26 , n28 , n29 , n30 , n31 , n34 , n36 , n38 , n40 , n43 , n45 , n46 , n47 , n49 , n51 , n52 , n53 , n54 , n56 , n57 , n58 , n60 , n61 , n63 , n64 , n65 , n67 , n69 , n70 , n71 , n72 , n73 , n74 , n76 , n77 , n78 , n79 , n80 , n81 , n83 , n84 , n85 , n86 , n87 , n90 , n93 , n94 , n95 , n97 , n99 , n103 , n105 , n106 , n108 , n109 , n111 , n112 , n113 , n114 , n116 , n117 , n118 , n120 , n121 , n122 , n123 , n125 , n127 , n128 , n129 , n130 , n131 , n133 , n135 , n137 , n139 , n140 , n141 , n143 , n144 , n145 , n146 , n148 , n151 , n152 , n153 , n155 , n157 , n158 , n160 , n161 , n163 , n164 , n165 , n167 , n168 , n169 , n171 , n173 , n174 , n175 , n176 , n178 , n180 , n182 , n184 , n185 , n186 , n187 , n189 , n191 , n192 , n194 , n195 , n198 , n199 , n200 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n210 , n211 , n212 , n213 , n214 , n216 , n217 , n218 , n219 , n221 , n222 , n223 , n225 , n227 , n228 , n231 , n232 , n235 , n236 , n238 , n241 , n242 , n243 , n244 , n245 , n247 , n248 , n249 , n252 , n253 , n255 , n256 , n258 , n259 , n260 , n261 , n262 , n263 , n265 , n267 , n268 , n271 , n272 , n273 , n275 , n276 , n277 , n278 , n280 , n282 , n283 , n285 , n286 , n287 , n288 , n290 , n291 , n292 , n293 , n295 , n296 , n297 , n299 , n300 , n301 , n303 , n304 , n306 , n307 , n308 , n310 , n312 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n334 , n335 , n336 , n337 , n338 , n339 , n341 , n342 , n343 , n344 , n346 , n347 , n348 , n349 , n351 , n352 , n353 , n354 , n356 , n357 , n358 , n360 , n361 , n362 , n363 , n364 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n374 , n375 , n376 , n377 , n378 , n380 , n382 , n383 , n384 , n386 , n387 , n388 , n389 , n391 , n392 , n396 , n397 , n398 , n399 , n401 , n402 , n403 , n404 , n406 , n407 , n408 , n409 , n410 , n411 , n413 , n415 , n416 , n418 , n419 , n421 , n425 , n426 , n427 , n429 , n430 , n432 , n434 , n436 , n437 , n439 , n440 , n442 , n443 , n444 , n445 , n447 , n448 , n450 , n451 , n453 , n455 , n457 , n459 , n462 , n463 , n464 , n465 , n466 , n468 , n469 , n471 , n473 , n474 , n475 , n476 , n478 , n479 , n481 , n482 , n484 , n485 , n486 , n488 , n489 , n490 , n492 , n493 , n495 , n496 , n497 , n498 , n501 , n502 , n503 , n505 , n507 , n508 , n510 , n511 , n512 , n513 , n516 , n518 , n519 , n521 , n522 , n523 , n524 , n525 , n527 , n529 , n530 , n532 , n533 , n534 , n537 , n538 , n539 , n541 , n542 , n544 , n546 , n549 , n551 , n552 , n554 , n556 , n558 , n559 , n561 , n563 , n564 , n565 , n566 , n570 , n571 , n572 , n573 , n575 , n576 , n578 , n580 , n581 , n583 , n584 , n585 , n586 , n589 , n590 , n591 , n593 , n594 , n595 , n596 , n598 , n600 , n602 , n604 , n605 , n606 , n607 , n608 , n610 , n611 , n613 , n614 , n615 , n619 , n620 , n621 , n622 , n624 , n626 , n628 , n629 , n630 , n632 , n636 , n638 , n639 , n640 , n641 , n642 , n644 , n645 , n647 , n648 , n650 , n651 , n652 , n654 , n656 , n657 , n658 , n660 , n661 , n662 , n665 , n667 , n669 , n671 , n672 , n674 , n676 , n678 , n681 , n682 , n684 , n685 , n686 , n690 , n692 , n694 , n695 , n697 , n698 , n700 , n701 , n703 , n705 , n706 , n707 , n709 , n710 , n713 , n714 , n716 , n718 , n719 , n721 , n724 , n727 , n730 , n732 , n733 , n734 , n736 , n737 , n738 , n740 , n741 , n742 , n743 , n744 , n746 , n747 , n748 , n750 , n751 , n752 , n753 , n754 , n756 , n757 , n758 , n759 , n761 , n762 , n763 , n765 , n770 , n771 , n772 , n773 , n774 , n776 , n777 , n778 , n780 , n781 , n782 , n784 , n787 , n788 , n790 , n791 , n792 , n794 , n795 , n797 , n798 , n800 , n801 , n802 , n805 , n806 , n808 , n809 , n810 , n812 , n813 , n815 , n817 , n818 , n819 , n824 , n825 , n826 , n827 , n830 , n833 , n835 , n836 , n838 , n839 , n841 , n842 , n844 , n846 , n847 , n848 , n851 , n854 , n856 , n858 , n860 , n861 , n863 , n864 , n865 , n866 , n868 , n869 , n870 , n872 , n874 , n875 , n876 , n878 , n879 , n880 , n883 , n886 , n889 , n890 , n891 , n895 , n896 , n897 , n899 , n900 , n902 , n903 , n905 , n906 , n908 , n910 , n911 , n913 , n914 , n916 , n917 , n918 , n919 , n921 , n922 , n923 , n925 , n926 , n929 , n930 , n931 , n934 , n935 , n936 , n938 , n939 , n940 , n943 , n945 , n947 , n948 , n949 , n950 , n951 , n953 , n955 , n957 , n959 , n961 , n962 , n963 , n964 , n965 , n967 , n968 , n969 , n970 , n971 , n972 , n974 , n975 , n976 , n977 , n978 , n980 , n981 , n982 , n983 , n984 , n987 , n988 , n989 , n990 , n993 , n994 , n995 , n997 , n998 , n999 , n1000 , n1001 , n1003 , n1004 , n1007 , n1008 , n1011 , n1012 , n1016 , n1017 , n1019 , n1020 , n1022 , n1023 , n1026 , n1027 , n1028 , n1029 , n1032 , n1033 , n1034 , n1036 , n1039 , n1040 , n1045 , n1046 , n1047 , n1050 , n1051 , n1054 , n1059 , n1060 , n1062 , n1064 , n1066 , n1068 , n1071 , n1075 , n1077 , n1078 , n1080 , n1082 , n1083 , n1087 , n1090 , n1092 , n1093 , n1095 , n1096 , n1102 , n1103 , n1106 , n1109 , n1110 , n1111 , n1112 , n1114 , n1115 , n1117 , n1118 , n1120 , n1121 , n1122 , n1125 , n1128 , n1132 , n1134 , n1135 , n1137 , n1138 , n1139 , n1140 , n1144 , n1145 , n1146 , n1150 , n1151 , n1154 , n1155 , n1158 , n1160 , n1161 , n1163 , n1164 , n1166 , n1167 , n1169 , n1173 , n1175 , n1176 , n1180 , n1182 , n1184 , n1186 , n1188 , n1189 , n1190 , n1191 , n1193 , n1195 , n1196 , n1197 , n1201 , n1203 , n1204 , n1205 , n1206 , n1208 , n1209 , n1210 , n1211 , n1213 , n1214 , n1215 , n1216 , n1218 , n1220 , n1222 , n1223 , n1226 , n1229 , n1231 , n1232 , n1234 , n1235 , n1237 , n1238 , n1240 , n1242 , n1245 , n1246 , n1247 , n1248 , n1250 , n1251 , n1253 , n1254 , n1255 , n1257 , n1258 , n1259 , n1261 , n1262 , n1263 , n1265 , n1266 , n1269 , n1271 , n1272 , n1275 , n1277 , n1278 , n1280 , n1283 , n1287 , n1289 , n1290 , n1291 , n1292 , n1294 , n1295 , n1296 , n1297 , n1299 , n1300 , n1301 , n1302 , n1303 , n1305 , n1306 , n1310 , n1311 , n1312 , n1314 , n1315 , n1317 , n1319 , n1320 , n1322 , n1324 , n1326 , n1329 , n1331 , n1332 , n1334 , n1336 , n1337 , n1339 , n1340 , n1342 , n1343 , n1345 , n1349 , n1352 , n1354 , n1356 , n1357 , n1358 , n1359 , n1361 , n1362 , n1363 , n1364 , n1370 , n1373 , n1376 , n1378 , n1380 , n1383 , n1385 , n1387 , n1389 , n1391 , n1393 , n1399 , n1400 , n1402 , n1403 , n1404 , n1405 , n1407 , n1408 , n1409 , n1410 , n1412 , n1414 , n1416 , n1419 , n1421 , n1422 , n1424 , n1426 , n1428 , n1429 , n1431 , n1432 , n1433 , n1434 , n1435 , n1437 , n1438 , n1440 , n1443 , n1445 , n1450 , n1451 , n1453 , n1454 , n1455 , n1457 , n1458 , n1460 , n1462 , n1463 , n1464 , n1466 , n1467 , n1469 , n1470 , n1471 , n1472 , n1475 , n1477 , n1478 , n1480 , n1482 , n1483 , n1484 , n1485 , n1489 , n1490 , n1492 , n1495 , n1496 , n1497 , n1499 , n1501 , n1502 , n1503 , n1505 , n1506 , n1509 , n1510 , n1511 , n1513 , n1514 , n1515 , n1517 , n1518 , n1521 , n1522 , n1525 , n1527 , n1528 , n1529 , n1530 , n1535 , n1536 , n1537 , n1540 , n1541 , n1542 , n1545 , n1546 , n1547 , n1549 , n1550 , n1551 , n1553 , n1554 , n1555 , n1556 , n1558 , n1559 , n1560 , n1562 , n1564 , n1565 , n1567 , n1568 , n1569 , n1570 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1579 , n1581 , n1582 , n1583 , n1584 , n1586 , n1587 , n1590 , n1594 , n1595 , n1596 , n1597 , n1598 , n1600 , n1601 , n1603 , n1604 , n1605 , n1606 , n1608 , n1610 , n1613 , n1614 , n1615 , n1617 , n1618 , n1619 , n1620 , n1623 , n1624 , n1625 , n1627 , n1629 , n1632 , n1635 , n1636 , n1637 , n1639 , n1640 , n1641 , n1643 , n1644 , n1646 , n1647 , n1649 , n1651 , n1653 , n1656 , n1657 , n1659 , n1660 , n1661 , n1664 , n1665 , n1667 , n1668 , n1669 , n1671 , n1672 , n1674 , n1675 , n1676 , n1678 , n1679 , n1680 , n1682 , n1683 , n1684 , n1685 , n1686 , n1688 , n1689 , n1690 , n1692 , n1693 , n1694 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1703 , n1704 , n1705 , n1707 , n1708 , n1712 , n1715 , n1717 , n1718 , n1720 , n1726 , n1727 , n1729 , n1730 , n1731 , n1737 , n1738 , n1739 , n1742 , n1743 , n1744 , n1745 , n1747 , n1748 , n1749 , n1750 , n1751 , n1755 , n1757 , n1758 , n1762 , n1766 , n1767 , n1768 , n1770 , n1772 , n1774 , n1775 , n1778 , n1779 , n1782 , n1785 , n1786 , n1787 , n1791 , n1793 , n1796 , n1798 , n1800 , n1802 , n1805 , n1809 , n1815 , n1817 , n1819 , n1825 , n1829 , n1830 , n1831 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1846 , n1851 , n1853 , n1858 , n1860 , n1862 , n1863 , n1870 , n1873 , n1874 , n1878 , n1879 , n1881 , n1885 , n1886 , n1887 , n1889 , n1891 , n1894 , n1896 , n1900 , n1903 , n1907 , n1910 , n1911 , n1912 , n1917 , n1920 , n1921 , n1923 , n1924 , n1927 , n1928 , n1932 , n1939 , n1942 , n1946 , n1948 , n1950 , n1952 , n1954 , n1956 , n1957 , n1959 , n1960 , n1963 , n1964 , n1967 , n1969 , n1970 , n1971 , n1974 , n1977 , n1980 , n1984 , n1989 , n1992 , n1995 , n1997 , n2001 , n2003 , n2005 , n2006 , n2008 , n2009 , n2013 , n2016 , n2017 , n2019 , n2020 , n2021 , n2022 , n2024 , n2025 , n2027 , n2028 , n2031 , n2036 , n2038 , n2040 , n2047 , n2049 , n2050 , n2051 , n2054 , n2059 , n2060 , n2063 , n2067 , n2068 , n2069 , n2070 , n2072 , n2073 , n2085 , n2090 , n2092 , n2095 , n2096 , n2097 , n2099 , n2104 , n2107 , n2113 , n2116 , n2117 , n2119 , n2121 , n2122 , n2123 , n2125 , n2126 , n2128 , n2131 , n2133 , n2134 , n2136 , n2137 , n2138 , n2140 , n2141 , n2145 , n2146 , n2147 , n2150 , n2154 , n2156 , n2158 , n2160 , n2162 , n2163 , n2164 , n2165 , n2169 , n2172 , n2173 , n2175 , n2176 , n2178 , n2180 , n2181 , n2182 , n2184 , n2189 , n2190 , n2193 , n2195 , n2199 , n2202 , n2204 , n2208 , n2210 , n2211 , n2212 , n2213 , n2215 , n2217 , n2218 , n2221 , n2222 , n2223 , n2224 , n2226 , n2227 , n2229 , n2231 , n2232 , n2235 , n2237 , n2239 , n2241 , n2242 , n2243 , n2245 , n2246 , n2249 , n2252 , n2254 , n2256 , n2258 , n2259 , n2261 , n2262 , n2263 , n2264 , n2265 , n2269 , n2271 , n2273 , n2274 , n2276 , n2277 , n2278 , n2279 , n2280 , n2282 , n2285 , n2287 , n2288 , n2291 , n2292 , n2294 , n2296 , n2298 , n2302 , n2306 , n2307 , n2309 , n2311 , n2312 , n2315 , n2317 , n2319 , n2321 , n2322 , n2323 , n2324 , n2326 , n2327 , n2328 , n2329 , n2331 , n2336 , n2338 , n2340 , n2341 , n2343 , n2345 , n2347 , n2351 , n2355 , n2356 , n2358 , n2359 , n2360 , n2362 , n2363 , n2364 , n2365 , n2366 , n2369 , n2370 , n2381 , n2383 , n2387 , n2391 , n2393 , n2394 , n2397 , n2398 , n2404 , n2405 , n2407 , n2410 , n2411 , n2412 , n2414 , n2415 , n2416 , n2418 , n2419 , n2421 , n2423 , n2424 , n2427 , n2432 , n2433 , n2434 , n2436 , n2437 , n2440 , n2441 , n2443 , n2445 , n2447 , n2449 , n2452 , n2454 , n2455 , n2456 , n2458 , n2462 , n2463 , n2465 , n2466 , n2467 , n2470 , n2471 , n2474 , n2475 , n2478 , n2479 , n2481 , n2489 , n2490 , n2493 , n2496 , n2498 , n2500 , n2503 , n2504 , n2507 , n2508 , n2509 , n2511 , n2513 , n2514 , n2516 , n2518 , n2522 , n2524 , n2527 , n2532 , n2534 , n2538 , n2540 , n2542 , n2544 , n2545 , n2546 , n2548 , n2549 , n2551 , n2552 , n2555 , n2556 , n2557 , n2559 , n2560 , n2562 , n2563 , n2565 , n2566 , n2567 , n2568 , n2569 , n2571 , n2572 , n2573 , n2575 , n2576 , n2577 , n2578 , n2579 , n2581 , n2583 , n2585 , n2587 , n2588 , n2590 , n2593 , n2594 , n2596 , n2597 , n2600 , n2602 , n2605 , n2607 , n2608 , n2610 , n2612 , n2619 , n2621 , n2623 , n2625 , n2629 , n2630 , n2639 , n2640 , n2641 , n2643 , n2645 , n2647 , n2650 , n2652 , n2657 , n2658 , n2661 , n2663 , n2665 , n2668 , n2672 , n2674 , n2675 , n2679 , n2684 , n2688 , n2693 , n2699 , n2701 , n2705 , n2706 , n2710 , n2711 , n2712 , n2714 , n2715 , n2716 , n2718 , n2719 , n2720 , n2721 , n2722 , n2724 , n2726 , n2728 , n2729 , n2731 , n2732 , n2734 , n2736 , n2738 , n2739 , n2740 , n2742 , n2743 , n2744 , n2746 , n2748 , n2749 , n2750 , n2752 , n2753 , n2754 , n2756 , n2757 , n2760 , n2761 , n2763 , n2765 , n2766 , n2767 , n2768 , n2772 , n2773 , n2775 , n2776 , n2777 , n2778 , n2779 , n2781 , n2782 , n2784 , n2785 , n2787 , n2788 , n2789 , n2790 , n2792 , n2793 , n2794 , n2796 , n2797 , n2800 , n2801 , n2802 , n2804 , n2807 , n2809 , n2810 , n2811 , n2813 , n2814 , n2818 , n2820 , n2825 , n2828 , n2830 , n2832 , n2833 , n2836 , n2839 , n2841 , n2843 , n2847 , n2848 , n2849 , n2853 , n2860 , n2865 , n2868 , n2871 , n2872 , n2873 , n2876 , n2877 , n2878 , n2879 , n2880 , n2882 , n2883 , n2885 , n2886 , n2887 , n2889 , n2891 , n2892 , n2893 , n2895 , n2896 , n2897 , n2898 , n2900 , n2902 , n2903 , n2904 , n2905 , n2906 , n2908 , n2910 , n2911 , n2913 , n2914 , n2915 , n2917 , n2918 , n2921 , n2922 , n2923 , n2924 , n2927 , n2931 , n2940 , n2948 , n2952 , n2953 , n2957 , n2959 , n2960 , n2963 , n2964 , n2965 , n2966 , n2969 , n2970 , n2971 , n2974 , n2977 , n2979 , n2980 , n2981 , n2982 , n2984 , n2986 , n2987 , n2989 , n2990 , n2992 , n2993 , n2994 , n2995 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3004 , n3005 , n3006 , n3007 , n3009 , n3011 , n3012 , n3013 , n3014 , n3016 , n3018 , n3019 , n3021 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3033 , n3034 , n3035 , n3036 , n3039 , n3040 , n3043 , n3045 , n3047 , n3049 , n3050 , n3054 , n3055 , n3057 , n3060 , n3061 , n3062 , n3064 , n3065 , n3069 , n3070 , n3072 , n3073 , n3077 , n3080 , n3083 , n3085 , n3089 , n3091 , n3093 , n3095 , n3097 , n3099 , n3101 , n3105 , n3107 , n3109 , n3112 , n3116 , n3117 , n3118 , n3119 , n3121 , n3123 , n3124 , n3128 , n3129 , n3132 , n3133 , n3134 , n3135 , n3138 , n3139 , n3141 , n3143 , n3144 , n3145 , n3147 , n3148 , n3149 , n3156 , n3157 , n3158 , n3160 , n3163 , n3164 , n3166 , n3168 , n3169 , n3170 , n3172 , n3173 , n3174 , n3176 , n3181 , n3182 , n3183 , n3184 , n3185 , n3189 , n3191 , n3192 , n3193 , n3195 , n3197 , n3198 , n3201 , n3203 , n3204 , n3207 , n3208 , n3209 , n3211 , n3212 , n3213 , n3215 , n3218 , n3222 , n3223 , n3224 , n3227 , n3228 , n3232 , n3234 , n3237 , n3238 , n3241 , n3243 , n3247 , n3249 , n3250 , n3251 , n3253 , n3256 , n3257 , n3259 , n3261 , n3263 , n3264 , n3265 , n3267 , n3268 , n3269 , n3271 , n3272 , n3274 , n3275 , n3276 , n3278 , n3279 , n3282 , n3284 , n3285 , n3286 , n3288 , n3290 , n3291 , n3292 , n3294 , n3295 , n3296 , n3297 , n3298 , n3301 , n3302 , n3304 , n3305 , n3307 , n3310 , n3311 , n3312 , n3315 , n3316 , n3317 , n3318 , n3321 , n3323 , n3325 , n3326 , n3327 , n3331 , n3333 , n3334 , n3336 , n3338 , n3341 , n3342 , n3344 , n3345 , n3349 , n3350 , n3354 , n3356 , n3359 , n3360 , n3361 , n3365 , n3366 , n3367 , n3369 , n3370 , n3371 , n3372 , n3374 , n3375 , n3376 , n3377 , n3380 , n3382 , n3384 , n3386 , n3387 , n3390 , n3391 , n3392 , n3394 , n3395 , n3398 , n3399 , n3404 , n3405 , n3406 , n3410 , n3412 , n3414 , n3415 , n3417 , n3423 , n3424 , n3426 , n3427 , n3428 , n3430 , n3433 , n3434 , n3436 , n3439 , n3443 , n3445 , n3446 , n3447 , n3448 , n3450 , n3453 , n3455 , n3457 , n3458 , n3459 , n3461 , n3462 , n3464 , n3466 , n3467 , n3469 , n3470 , n3471 , n3472 , n3474 , n3475 , n3476 , n3477 , n3478 , n3480 , n3482 , n3485 , n3486 , n3487 , n3488 , n3490 , n3491 , n3492 , n3493 , n3494 , n3496 , n3497 , n3498 , n3502 , n3504 , n3508 , n3509 , n3511 , n3512 , n3513 , n3515 , n3519 , n3520 , n3521 , n3523 , n3524 , n3525 , n3526 , n3527 , n3529 , n3536 , n3539 , n3541 , n3542 , n3548 , n3549 , n3550 , n3552 , n3556 , n3558 , n3561 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3570 , n3571 , n3572 , n3574 , n3576 , n3577 , n3579 , n3580 , n3581 , n3584 , n3585 , n3586 , n3588 , n3589 , n3590 , n3592 , n3594 , n3595 , n3598 , n3599 , n3600 , n3601 , n3603 , n3604 , n3605 , n3606 , n3608 , n3609 , n3611 , n3612 , n3613 , n3617 , n3618 , n3620 , n3621 , n3622 , n3624 , n3625 , n3626 , n3628 , n3629 , n3630 , n3632 , n3634 , n3636 , n3637 , n3638 , n3640 , n3641 , n3642 , n3645 , n3646 , n3647 , n3648 , n3649 , n3652 , n3655 , n3657 , n3659 , n3660 , n3661 , n3662 , n3666 , n3667 , n3677 , n3678 , n3681 , n3683 , n3685 , n3687 , n3688 , n3692 , n3694 , n3696 , n3700 , n3701 , n3702 , n3703 , n3705 , n3706 , n3710 , n3712 , n3713 , n3715 , n3718 , n3719 , n3721 , n3723 , n3724 , n3726 , n3732 , n3736 , n3738 , n3739 , n3741 , n3742 , n3744 , n3747 , n3748 , n3750 , n3751 , n3754 , n3755 , n3761 , n3762 , n3763 , n3766 , n3774 , n3776 , n3777 , n3778 , n3780 , n3781 , n3784 , n3785 , n3786 , n3789 , n3790 , n3792 , n3794 , n3796 , n3797 , n3799 , n3800 , n3802 , n3804 , n3805 , n3807 , n3808 , n3810 , n3811 , n3817 , n3818 , n3819 , n3820 , n3823 , n3824 , n3825 , n3826 , n3828 , n3829 , n3830 , n3832 , n3833 , n3834 , n3835 , n3837 , n3840 , n3841 , n3842 , n3843 , n3845 , n3847 , n3848 , n3850 , n3852 , n3854 , n3855 , n3857 , n3859 , n3860 , n3862 , n3863 , n3864 , n3866 , n3867 , n3871 , n3874 , n3879 , n3880 , n3882 , n3883 , n3884 , n3890 , n3891 , n3892 , n3893 , n3896 , n3897 , n3898 , n3899 , n3901 , n3902 , n3903 , n3905 , n3906 , n3907 , n3909 , n3914 , n3918 , n3919 , n3922 , n3924 , n3927 , n3929 , n3930 , n3934 , n3936 , n3937 , n3939 , n3940 , n3943 , n3944 , n3946 , n3948 , n3949 , n3951 , n3955 , n3960 , n3963 , n3965 , n3966 , n3968 , n3971 , n3974 , n3977 , n3978 , n3979 , n3981 , n3983 , n3984 , n3987 , n3989 , n3990 , n3992 , n3993 , n3997 , n3999 , n4000 , n4005 , n4006 , n4009 , n4010 , n4011 , n4014 , n4015 , n4016 , n4018 , n4019 , n4022 , n4024 , n4026 , n4028 , n4030 , n4031 , n4033 , n4034 , n4035 , n4037 , n4038 , n4039 , n4042 , n4047 , n4048 , n4050 , n4052 , n4055 , n4056 , n4057 , n4059 , n4061 , n4062 , n4065 , n4068 , n4070 , n4075 , n4076 , n4077 , n4078 , n4081 , n4082 , n4083 , n4085 , n4086 , n4088 , n4089 , n4090 , n4094 , n4096 , n4099 , n4100 , n4101 , n4102 , n4103 , n4105 , n4107 , n4108 , n4109 , n4111 , n4114 , n4116 , n4117 , n4118 , n4122 , n4124 , n4129 , n4130 , n4131 , n4136 , n4137 , n4139 , n4142 , n4149 , n4150 , n4151 , n4155 , n4162 , n4165 , n4166 , n4167 , n4171 , n4173 , n4175 , n4180 , n4188 , n4189 , n4190 , n4192 , n4195 , n4197 , n4200 , n4201 , n4202 , n4203 , n4205 , n4209 , n4211 , n4212 , n4213 , n4216 , n4217 , n4219 , n4225 , n4228 , n4230 , n4232 , n4233 , n4234 , n4235 , n4238 , n4239 , n4240 , n4241 , n4243 , n4246 , n4249 , n4250 , n4253 , n4254 , n4259 , n4260 , n4261 , n4262 , n4263 , n4265 , n4269 , n4270 , n4273 , n4274 , n4275 , n4276 , n4279 , n4280 , n4282 , n4285 , n4286 , n4288 , n4289 , n4291 , n4293 , n4294 , n4295 , n4298 , n4299 , n4300 , n4302 , n4304 , n4305 , n4306 , n4308 , n4312 , n4313 , n4314 , n4317 , n4320 , n4321 , n4325 , n4326 , n4329 , n4331 , n4335 , n4336 , n4338 , n4340 , n4341 , n4349 , n4351 , n4353 , n4357 , n4360 , n4361 , n4362 , n4366 , n4368 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4380 , n4382 , n4383 , n4387 , n4389 , n4392 , n4395 , n4399 , n4401 , n4403 , n4409 , n4411 , n4412 , n4415 , n4416 , n4417 , n4419 , n4420 , n4422 , n4423 , n4424 , n4426 , n4429 , n4431 , n4432 , n4433 , n4438 , n4439 , n4441 , n4443 , n4444 , n4448 , n4451 , n4453 , n4455 , n4457 , n4459 , n4460 , n4463 , n4465 , n4467 , n4469 , n4475 , n4478 , n4479 , n4482 , n4483 , n4486 , n4487 , n4489 , n4490 , n4494 , n4495 , n4497 , n4502 , n4504 , n4507 , n4508 , n4514 , n4515 , n4518 , n4519 , n4520 , n4523 , n4526 , n4527 , n4528 , n4529 , n4532 , n4535 , n4536 , n4540 , n4541 , n4543 , n4545 , n4548 , n4550 , n4551 , n4552 , n4554 , n4559 , n4561 , n4562 , n4564 , n4567 , n4569 , n4570 , n4571 , n4572 , n4573 , n4575 , n4576 , n4581 , n4583 , n4584 , n4586 , n4587 , n4588 , n4589 , n4591 , n4594 , n4595 , n4596 , n4598 , n4601 , n4602 , n4604 , n4606 , n4607 , n4608 , n4611 , n4612 , n4614 , n4615 , n4618 , n4619 , n4621 , n4625 , n4626 , n4627 , n4631 , n4632 , n4633 , n4635 , n4636 , n4638 , n4640 , n4643 , n4644 , n4647 , n4648 , n4649 , n4651 , n4654 , n4656 , n4657 , n4660 , n4662 , n4665 , n4666 , n4667 , n4668 , n4670 , n4672 , n4674 , n4678 , n4679 , n4681 , n4683 , n4684 , n4688 , n4689 , n4693 , n4695 , n4699 , n4702 , n4703 , n4708 , n4709 , n4714 , n4719 , n4720 , n4723 , n4726 , n4727 , n4728 , n4731 , n4732 , n4734 , n4736 , n4737 , n4739 , n4740 , n4745 , n4748 , n4751 , n4753 , n4754 , n4755 , n4757 , n4758 , n4763 , n4764 , n4765 , n4766 , n4768 , n4771 , n4775 , n4777 , n4780 , n4781 , n4784 , n4788 , n4789 , n4792 , n4795 , n4804 , n4808 , n4811 , n4815 , n4816 , n4817 , n4818 , n4820 , n4821 , n4822 , n4824 , n4828 , n4830 , n4831 , n4833 , n4835 , n4840 , n4841 , n4843 , n4844 , n4847 , n4849 , n4850 , n4853 , n4855 , n4856 , n4861 , n4864 , n4868 , n4874 , n4876 , n4877 , n4878 , n4882 , n4885 , n4889 , n4891 , n4892 , n4895 , n4898 , n4903 , n4904 , n4907 , n4908 , n4910 , n4911 , n4914 , n4915 , n4916 , n4917 , n4918 , n4920 , n4921 , n4922 , n4924 , n4925 , n4926 , n4931 , n4932 , n4933 , n4935 , n4937 , n4938 , n4940 , n4942 , n4945 , n4948 , n4949 , n4950 , n4951 , n4953 , n4954 , n4957 , n4959 , n4960 , n4961 , n4962 , n4964 , n4972 , n4973 , n4976 , n4977 , n4978 , n4979 , n4981 , n4982 , n4983 , n4987 , n4990 , n4991 , n4995 , n4998 , n5001 , n5003 , n5004 , n5007 , n5008 , n5009 , n5012 , n5014 , n5016 , n5017 , n5022 , n5030 , n5032 , n5033 , n5034 , n5035 , n5037 , n5039 , n5040 , n5048 , n5049 , n5054 , n5055 , n5056 , n5057 , n5059 , n5061 , n5064 , n5065 , n5066 , n5072 , n5076 , n5077 , n5080 , n5081 , n5084 , n5085 , n5086 , n5087 , n5088 , n5090 , n5091 , n5094 , n5095 , n5097 , n5098 , n5099 , n5101 , n5103 , n5105 , n5106 , n5108 , n5109 , n5111 , n5114 , n5116 , n5117 , n5120 , n5124 , n5125 , n5127 , n5128 , n5129 , n5132 , n5140 , n5141 , n5143 , n5145 , n5148 , n5151 , n5153 , n5159 , n5161 , n5164 , n5166 , n5167 , n5173 , n5174 , n5176 , n5177 , n5178 , n5179 , n5181 , n5183 , n5184 , n5186 , n5190 , n5193 , n5201 , n5209 , n5210 , n5212 , n5213 , n5214 , n5215 , n5217 , n5224 , n5227 , n5228 , n5229 , n5233 , n5235 , n5236 , n5237 , n5239 , n5243 , n5244 , n5245 , n5247 , n5250 , n5251 , n5253 , n5256 , n5257 , n5259 , n5261 , n5266 , n5269 , n5270 , n5271 , n5273 , n5274 , n5278 , n5279 , n5281 , n5285 , n5286 , n5288 , n5293 , n5294 , n5296 , n5297 , n5303 , n5304 , n5305 , n5307 , n5310 , n5314 , n5318 , n5320 , n5323 , n5324 , n5326 , n5329 , n5331 , n5333 , n5335 , n5337 , n5342 , n5345 , n5349 , n5351 , n5354 , n5355 , n5357 , n5362 , n5363 , n5366 , n5368 , n5370 , n5372 , n5373 , n5378 , n5380 , n5381 , n5382 , n5385 , n5390 , n5393 , n5398 , n5399 , n5401 , n5403 , n5410 , n5411 , n5413 , n5417 , n5419 , n5422 , n5423 , n5424 , n5425 , n5427 , n5433 , n5435 , n5438 , n5440 , n5441 , n5442 , n5443 , n5446 , n5449 , n5451 , n5457 , n5461 , n5463 , n5465 , n5466 , n5471 , n5476 , n5477 , n5479 , n5482 , n5483 , n5484 , n5493 , n5495 , n5497 , n5499 , n5507 , n5510 , n5513 , n5514 , n5516 , n5518 , n5520 , n5522 , n5529 , n5531 , n5534 , n5536 , n5539 , n5543 , n5544 , n5547 , n5550 , n5553 , n5554 , n5557 , n5558 , n5564 , n5565 , n5568 , n5569 , n5574 , n5575 , n5586 , n5587 , n5589 , n5595 , n5598 , n5603 , n5606 , n5609 , n5611 , n5613 , n5619 , n5628 , n5630 , n5631 , n5633 , n5636 , n5637 , n5640 , n5641 , n5643 , n5647 , n5650 , n5651 , n5652 , n5654 , n5661 , n5665 , n5666 , n5667 , n5670 , n5673 , n5677 , n5678 , n5679 , n5680 , n5681 , n5683 , n5686 , n5688 , n5689 , n5690 , n5692 , n5693 , n5696 , n5697 , n5700 , n5701 , n5703 , n5704 , n5707 , n5711 , n5716 , n5718 , n5720 , n5727 , n5730 , n5732 , n5733 , n5734 , n5735 , n5736 , n5738 , n5739 , n5740 , n5744 , n5752 , n5754 , n5756 , n5758 , n5759 , n5763 , n5764 , n5766 , n5767 , n5768 , n5770 , n5773 , n5775 , n5776 , n5777 , n5779 , n5790 , n5798 , n5800 , n5801 , n5802 , n5808 , n5809 , n5811 , n5812 , n5816 , n5819 , n5825 , n5827 , n5828 , n5830 , n5832 , n5833 , n5839 , n5840 , n5841 , n5843 , n5853 , n5854 , n5855 , n5857 , n5858 , n5859 , n5862 , n5867 , n5868 , n5869 , n5870 , n5876 , n5877 , n5879 , n5884 , n5886 , n5889 , n5892 , n5893 , n5894 , n5903 , n5904 , n5905 , n5906 , n5910 , n5916 , n5918 , n5926 , n5928 , n5929 , n5931 , n5932 , n5939 , n5941 , n5942 , n5951 , n5952 , n5956 , n5957 , n5963 , n5964 , n5968 , n5969 , n5972 , n5976 , n5978 , n5980 , n5981 , n5985 , n5987 , n5990 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n6000 , n6001 , n6004 , n6010 , n6011 , n6014 , n6019 , n6025 , n6033 , n6035 , n6036 , n6040 , n6041 , n6043 , n6045 , n6048 , n6060 , n6061 , n6064 , n6065 , n6066 , n6067 , n6068 , n6073 , n6079 , n6080 , n6085 , n6087 , n6091 , n6097 , n6103 , n6105 , n6107 , n6108 , n6109 , n6112 , n6115 , n6116 , n6118 , n6119 , n6122 , n6123 , n6125 , n6126 , n6128 , n6131 , n6134 , n6137 , n6138 , n6139 , n6141 , n6150 , n6151 , n6157 , n6158 , n6159 , n6160 , n6162 , n6163 , n6170 , n6173 , n6174 , n6176 , n6177 , n6185 , n6186 , n6187 , n6190 , n6192 , n6196 , n6198 , n6199 , n6202 , n6204 , n6206 , n6212 , n6218 , n6220 , n6223 , n6228 , n6229 , n6230 , n6233 , n6234 , n6235 , n6236 , n6237 , n6239 , n6240 , n6241 , n6245 , n6247 , n6249 , n6252 , n6253 , n6254 , n6256 , n6258 , n6259 , n6260 , n6264 , n6265 , n6266 , n6269 , n6271 , n6272 , n6274 , n6275 , n6277 , n6278 , n6282 , n6285 , n6287 , n6291 , n6292 , n6293 , n6295 , n6301 , n6304 , n6306 , n6307 , n6308 , n6310 , n6313 , n6315 , n6322 , n6323 , n6326 , n6329 , n6331 , n6332 , n6334 , n6336 , n6337 , n6340 , n6341 , n6343 , n6344 , n6348 , n6349 , n6351 , n6357 , n6359 , n6360 , n6365 , n6367 , n6368 , n6371 , n6372 , n6373 , n6375 , n6378 , n6379 , n6382 , n6385 , n6387 , n6390 , n6393 , n6396 , n6398 , n6401 , n6403 , n6404 , n6405 , n6407 , n6413 , n6415 , n6418 , n6420 , n6422 , n6425 , n6426 , n6427 , n6429 , n6434 , n6435 , n6436 , n6437 , n6438 , n6441 , n6443 , n6446 , n6449 , n6452 , n6454 , n6455 , n6456 , n6460 , n6461 , n6463 , n6466 , n6469 , n6472 , n6473 , n6476 , n6480 , n6482 , n6487 , n6489 , n6492 , n6495 , n6497 , n6500 , n6504 , n6511 , n6515 , n6517 , n6520 , n6522 , n6524 , n6525 , n6528 , n6534 , n6535 , n6536 , n6539 , n6542 , n6545 , n6548 , n6551 , n6556 , n6558 , n6560 , n6563 , n6566 , n6569 , n6572 , n6576 , n6579 , n6582 , n6584 , n6586 , n6591 , n6592 , n6593 , n6594 , n6595 , n6601 , n6604 , n6606 , n6607 , n6609 , n6610 , n6612 , n6613 , n6615 , n6617 , n6624 , n6634 , n6635 , n6643 , n6645 , n6647 , n6651 , n6654 , n6657 , n6659 , n6664 , n6666 , n6667 , n6675 , n6678 , n6679 , n6682 , n6683 , n6687 , n6689 , n6690 , n6693 , n6694 , n6696 , n6698 , n6701 , n6703 , n6709 , n6713 , n6715 , n6719 , n6727 , n6729 , n6730 , n6731 , n6733 , n6737 , n6739 , n6746 , n6747 , n6748 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6774 , n6775 , n6776 , n6778 , n6779 , n6782 , n6783 , n6784 , n6787 , n6792 , n6798 , n6802 , n6803 , n6808 , n6809 , n6810 , n6814 , n6815 , n6818 , n6819 , n6821 , n6825 , n6831 , n6832 , n6834 , n6837 , n6839 , n6840 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6851 , n6856 , n6858 , n6860 , n6863 , n6865 , n6866 , n6867 , n6868 , n6870 , n6871 , n6873 , n6876 , n6877 , n6881 , n6882 , n6884 , n6887 , n6888 , n6890 , n6891 , n6892 , n6894 , n6897 , n6900 , n6902 , n6903 , n6905 , n6906 , n6908 , n6909 , n6910 , n6912 , n6914 , n6915 , n6926 , n6928 , n6931 , n6933 , n6934 , n6936 , n6941 , n6944 , n6952 , n6953 , n6958 , n6960 , n6964 , n6966 , n6970 , n6971 , n6972 , n6975 , n6977 , n6978 , n6983 , n6985 , n6988 , n6989 , n6991 , n6994 , n6999 , n7001 , n7010 , n7013 , n7015 , n7017 , n7019 , n7025 , n7026 , n7030 , n7033 , n7037 , n7038 , n7039 , n7040 , n7042 , n7044 , n7046 , n7048 , n7053 , n7054 , n7055 , n7056 , n7060 , n7063 , n7067 , n7074 , n7085 , n7099 , n7107 , n7108 , n7109 , n7114 , n7117 , n7122 , n7126 , n7129 , n7130 , n7131 , n7133 , n7134 , n7135 , n7137 , n7144 , n7145 , n7146 , n7148 , n7152 , n7155 , n7159 , n7162 , n7167 , n7168 , n7172 , n7182 , n7185 , n7188 , n7194 , n7196 , n7197 , n7198 , n7202 , n7205 , n7207 , n7209 , n7211 , n7214 , n7216 , n7218 , n7224 , n7225 , n7226 , n7229 , n7232 , n7235 , n7236 , n7237 , n7240 , n7241 , n7247 , n7249 , n7257 , n7260 , n7263 , n7265 , n7267 , n7273 , n7274 , n7276 , n7278 , n7282 , n7283 , n7290 , n7292 , n7293 , n7295 , n7297 , n7299 , n7306 , n7307 , n7314 , n7320 , n7322 , n7324 , n7326 , n7328 , n7331 , n7336 , n7338 , n7339 , n7343 , n7346 , n7350 , n7352 , n7355 , n7361 , n7362 , n7374 , n7375 , n7378 , n7380 , n7383 , n7392 , n7395 , n7397 , n7399 , n7403 , n7406 , n7409 , n7411 , n7412 , n7414 , n7415 , n7416 , n7418 , n7421 , n7422 , n7423 , n7427 , n7428 , n7430 , n7432 , n7433 , n7435 , n7438 , n7442 , n7444 , n7447 , n7448 , n7449 , n7451 , n7454 , n7455 , n7457 , n7461 , n7467 , n7468 , n7470 , n7474 , n7479 , n7481 , n7483 , n7484 , n7485 , n7486 , n7488 , n7489 , n7490 , n7494 , n7500 , n7501 , n7505 , n7506 , n7509 , n7514 , n7516 , n7519 , n7521 , n7523 , n7524 , n7526 , n7527 , n7528 , n7529 , n7532 , n7533 , n7535 , n7536 , n7537 , n7539 , n7543 , n7544 , n7545 , n7547 , n7548 , n7549 , n7551 , n7554 , n7556 , n7561 , n7562 , n7565 , n7566 , n7568 , n7571 , n7574 , n7581 , n7582 , n7585 , n7588 , n7589 , n7590 , n7591 , n7593 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7603 , n7604 , n7605 , n7609 , n7611 , n7615 , n7617 , n7619 , n7621 , n7623 , n7625 , n7627 , n7628 , n7631 , n7633 , n7637 , n7642 , n7644 , n7645 , n7648 , n7649 , n7650 , n7651 , n7653 , n7654 , n7656 , n7658 , n7660 , n7664 , n7665 , n7669 , n7673 , n7674 , n7675 , n7679 , n7681 , n7684 , n7687 , n7692 , n7694 , n7698 , n7704 , n7705 , n7708 , n7709 , n7710 , n7712 , n7716 , n7718 , n7719 , n7722 , n7728 , n7730 , n7739 , n7742 , n7747 , n7748 , n7751 , n7752 , n7756 , n7757 , n7758 , n7761 , n7763 , n7767 ;
  OR3x1_ASAP7_75t_R    g0000( .A (x2), .B (x1), .C (x0), .Y (y0) );
  AO21x1_ASAP7_75t_R   g0001( .A1 (x3), .A2 (x2), .B (x0), .Y (n9) );
  NOR2x1_ASAP7_75t_R   g0002( .A (x1), .B (n9), .Y (n10) );
  INVx1_ASAP7_75t_R    g0003( .A (n10), .Y (y1) );
  INVx1_ASAP7_75t_R    g0004( .A (x0), .Y (n12) );
  AND2x2_ASAP7_75t_R   g0005( .A (x2), .B (x1), .Y (n13) );
  INVx1_ASAP7_75t_R    g0006( .A (n13), .Y (n14) );
  INVx1_ASAP7_75t_R    g0007( .A (x2), .Y (n15) );
  INVx1_ASAP7_75t_R    g0008( .A (x1), .Y (n16) );
  INVx1_ASAP7_75t_R    g0009( .A (x3), .Y (n17) );
  AO21x1_ASAP7_75t_R   g0010( .A1 (n15), .A2 (n16), .B (n17), .Y (n18) );
  OR3x1_ASAP7_75t_R    g0011( .A (x2), .B (x1), .C (x3), .Y (n19) );
  AND3x1_ASAP7_75t_R   g0012( .A (n14), .B (n18), .C (n19), .Y (n20) );
  NAND2x1_ASAP7_75t_R  g0013( .A (n12), .B (n20), .Y (y2) );
  INVx1_ASAP7_75t_R    g0014( .A (x4), .Y (n22) );
  AO21x1_ASAP7_75t_R   g0015( .A1 (n22), .A2 (x5), .B (x0), .Y (n23) );
  INVx1_ASAP7_75t_R    g0016( .A (x5), .Y (y2079) );
  AO21x1_ASAP7_75t_R   g0017( .A1 (y2079), .A2 (x4), .B (x1), .Y (n25) );
  NOR2x1_ASAP7_75t_R   g0018( .A (n23), .B (n25), .Y (n26) );
  INVx1_ASAP7_75t_R    g0019( .A (n26), .Y (y3) );
  NAND2x1_ASAP7_75t_R  g0020( .A (x5), .B (n22), .Y (n28) );
  INVx1_ASAP7_75t_R    g0021( .A (n28), .Y (n29) );
  AO21x1_ASAP7_75t_R   g0022( .A1 (n16), .A2 (x5), .B (n22), .Y (n30) );
  INVx1_ASAP7_75t_R    g0023( .A (n30), .Y (n31) );
  OR3x1_ASAP7_75t_R    g0024( .A (n29), .B (n31), .C (x0), .Y (y4) );
  AND2x2_ASAP7_75t_R   g0025( .A (x1), .B (x0), .Y (y863) );
  AO21x1_ASAP7_75t_R   g0026( .A1 (x4), .A2 (x5), .B (y863), .Y (n34) );
  NOR2x1_ASAP7_75t_R   g0027( .A (x4), .B (x5), .Y (y2466) );
  AO21x1_ASAP7_75t_R   g0028( .A1 (n16), .A2 (n12), .B (y2466), .Y (n36) );
  NAND2x1_ASAP7_75t_R  g0029( .A (n34), .B (n36), .Y (y5) );
  AND3x1_ASAP7_75t_R   g0030( .A (n16), .B (n12), .C (x5), .Y (n38) );
  INVx1_ASAP7_75t_R    g0031( .A (n38), .Y (y6) );
  OR3x1_ASAP7_75t_R    g0032( .A (y863), .B (x5), .C (x2), .Y (n40) );
  AND2x2_ASAP7_75t_R   g0033( .A (n40), .B (y6), .Y (y7) );
  OR3x1_ASAP7_75t_R    g0034( .A (y2466), .B (x1), .C (x0), .Y (y8) );
  NOR2x1_ASAP7_75t_R   g0035( .A (x0), .B (x1), .Y (n43) );
  INVx1_ASAP7_75t_R    g0036( .A (n43), .Y (y9) );
  NOR2x1_ASAP7_75t_R   g0037( .A (x2), .B (x3), .Y (n45) );
  OR3x1_ASAP7_75t_R    g0038( .A (n45), .B (x1), .C (x0), .Y (n46) );
  OR3x1_ASAP7_75t_R    g0039( .A (n43), .B (x3), .C (x2), .Y (n47) );
  AND2x2_ASAP7_75t_R   g0040( .A (n46), .B (n47), .Y (y10) );
  AO21x1_ASAP7_75t_R   g0041( .A1 (n16), .A2 (n12), .B (n45), .Y (n49) );
  INVx1_ASAP7_75t_R    g0042( .A (n49), .Y (y11) );
  NOR2x1_ASAP7_75t_R   g0043( .A (x2), .B (x1), .Y (n51) );
  INVx1_ASAP7_75t_R    g0044( .A (n51), .Y (n52) );
  AND3x1_ASAP7_75t_R   g0045( .A (n15), .B (n16), .C (x5), .Y (n53) );
  AO21x1_ASAP7_75t_R   g0046( .A1 (y2079), .A2 (n52), .B (n53), .Y (n54) );
  OR3x1_ASAP7_75t_R    g0047( .A (n54), .B (n13), .C (x0), .Y (y12) );
  AO21x1_ASAP7_75t_R   g0048( .A1 (n12), .A2 (n16), .B (n15), .Y (n56) );
  INVx1_ASAP7_75t_R    g0049( .A (n56), .Y (n57) );
  AND2x2_ASAP7_75t_R   g0050( .A (x0), .B (x5), .Y (n58) );
  AO21x1_ASAP7_75t_R   g0051( .A1 (y2079), .A2 (x1), .B (n58), .Y (y2389) );
  OR3x1_ASAP7_75t_R    g0052( .A (x0), .B (x1), .C (x2), .Y (n60) );
  INVx1_ASAP7_75t_R    g0053( .A (n60), .Y (n61) );
  OR3x1_ASAP7_75t_R    g0054( .A (n57), .B (y2389), .C (n61), .Y (y13) );
  NAND2x1_ASAP7_75t_R  g0055( .A (x1), .B (n15), .Y (n63) );
  NAND2x1_ASAP7_75t_R  g0056( .A (x2), .B (n16), .Y (n64) );
  AND3x1_ASAP7_75t_R   g0057( .A (n63), .B (n64), .C (n12), .Y (n65) );
  AO21x1_ASAP7_75t_R   g0058( .A1 (n19), .A2 (x0), .B (n65), .Y (y14) );
  AO21x1_ASAP7_75t_R   g0059( .A1 (n15), .A2 (n16), .B (x0), .Y (n67) );
  AO21x1_ASAP7_75t_R   g0060( .A1 (n67), .A2 (n19), .B (n13), .Y (y15) );
  AO21x1_ASAP7_75t_R   g0061( .A1 (n17), .A2 (x2), .B (x0), .Y (n69) );
  AND3x1_ASAP7_75t_R   g0062( .A (n17), .B (x2), .C (x0), .Y (n70) );
  INVx1_ASAP7_75t_R    g0063( .A (n70), .Y (n71) );
  NAND2x1_ASAP7_75t_R  g0064( .A (x3), .B (n15), .Y (n72) );
  AND3x1_ASAP7_75t_R   g0065( .A (n16), .B (n15), .C (x3), .Y (n73) );
  AO21x1_ASAP7_75t_R   g0066( .A1 (n72), .A2 (x1), .B (n73), .Y (n74) );
  AO21x1_ASAP7_75t_R   g0067( .A1 (n69), .A2 (n71), .B (n74), .Y (y16) );
  AND2x2_ASAP7_75t_R   g0068( .A (x3), .B (x2), .Y (n76) );
  INVx1_ASAP7_75t_R    g0069( .A (n76), .Y (n77) );
  AND3x1_ASAP7_75t_R   g0070( .A (n16), .B (x2), .C (x3), .Y (n78) );
  AO21x1_ASAP7_75t_R   g0071( .A1 (n77), .A2 (x1), .B (n78), .Y (n79) );
  INVx1_ASAP7_75t_R    g0072( .A (n79), .Y (n80) );
  NOR2x1_ASAP7_75t_R   g0073( .A (x3), .B (x2), .Y (n81) );
  OR3x1_ASAP7_75t_R    g0074( .A (n80), .B (n81), .C (x0), .Y (y17) );
  AND2x2_ASAP7_75t_R   g0075( .A (n64), .B (n63), .Y (n83) );
  NAND2x1_ASAP7_75t_R  g0076( .A (x3), .B (n12), .Y (n84) );
  AND3x1_ASAP7_75t_R   g0077( .A (n12), .B (x2), .C (x1), .Y (n85) );
  INVx1_ASAP7_75t_R    g0078( .A (n85), .Y (n86) );
  AO21x1_ASAP7_75t_R   g0079( .A1 (n86), .A2 (n52), .B (x3), .Y (n87) );
  OA21x2_ASAP7_75t_R   g0080( .A1 (n83), .A2 (n84), .B (n87), .Y (y18) );
  OR3x1_ASAP7_75t_R    g0081( .A (n13), .B (y2079), .C (x0), .Y (y19) );
  NAND2x1_ASAP7_75t_R  g0082( .A (x0), .B (n16), .Y (n90) );
  AO21x1_ASAP7_75t_R   g0083( .A1 (n90), .A2 (y2079), .B (n58), .Y (y199) );
  AO21x1_ASAP7_75t_R   g0084( .A1 (x2), .A2 (y9), .B (y199), .Y (y20) );
  OR3x1_ASAP7_75t_R    g0085( .A (x2), .B (x1), .C (x5), .Y (n93) );
  INVx1_ASAP7_75t_R    g0086( .A (n93), .Y (n94) );
  INVx1_ASAP7_75t_R    g0087( .A (y19), .Y (n95) );
  NOR2x1_ASAP7_75t_R   g0088( .A (n94), .B (n95), .Y (y21) );
  NAND2x1_ASAP7_75t_R  g0089( .A (x5), .B (n15), .Y (n97) );
  AO21x1_ASAP7_75t_R   g0090( .A1 (n97), .A2 (n64), .B (x0), .Y (y22) );
  AO21x1_ASAP7_75t_R   g0091( .A1 (n15), .A2 (x5), .B (n16), .Y (n99) );
  NAND2x1_ASAP7_75t_R  g0092( .A (n12), .B (n99), .Y (y23) );
  OR3x1_ASAP7_75t_R    g0093( .A (n94), .B (n13), .C (x0), .Y (y24) );
  AO21x1_ASAP7_75t_R   g0094( .A1 (x2), .A2 (x1), .B (x0), .Y (y25) );
  AND2x2_ASAP7_75t_R   g0095( .A (x1), .B (x2), .Y (n103) );
  AO21x1_ASAP7_75t_R   g0096( .A1 (n71), .A2 (n84), .B (n103), .Y (y26) );
  AO21x1_ASAP7_75t_R   g0097( .A1 (n15), .A2 (x3), .B (n16), .Y (n105) );
  INVx1_ASAP7_75t_R    g0098( .A (n105), .Y (n106) );
  AO21x1_ASAP7_75t_R   g0099( .A1 (n71), .A2 (n69), .B (n106), .Y (y27) );
  OR3x1_ASAP7_75t_R    g0100( .A (x0), .B (x2), .C (x1), .Y (n108) );
  INVx1_ASAP7_75t_R    g0101( .A (n108), .Y (n109) );
  AO21x1_ASAP7_75t_R   g0102( .A1 (y19), .A2 (n93), .B (n109), .Y (y28) );
  NOR2x1_ASAP7_75t_R   g0103( .A (x1), .B (x3), .Y (n111) );
  INVx1_ASAP7_75t_R    g0104( .A (n111), .Y (n112) );
  AO21x1_ASAP7_75t_R   g0105( .A1 (x1), .A2 (x2), .B (x0), .Y (n113) );
  NOR2x1_ASAP7_75t_R   g0106( .A (x3), .B (n113), .Y (n114) );
  AO21x1_ASAP7_75t_R   g0107( .A1 (n112), .A2 (n113), .B (n114), .Y (y29) );
  AO21x1_ASAP7_75t_R   g0108( .A1 (n16), .A2 (n17), .B (x0), .Y (n116) );
  AND3x1_ASAP7_75t_R   g0109( .A (n16), .B (n17), .C (x2), .Y (n117) );
  NAND2x1_ASAP7_75t_R  g0110( .A (x0), .B (n117), .Y (n118) );
  OA21x2_ASAP7_75t_R   g0111( .A1 (n103), .A2 (n116), .B (n118), .Y (y30) );
  AO21x1_ASAP7_75t_R   g0112( .A1 (n16), .A2 (x3), .B (n15), .Y (n120) );
  NAND2x1_ASAP7_75t_R  g0113( .A (n12), .B (n120), .Y (n121) );
  AND3x1_ASAP7_75t_R   g0114( .A (n16), .B (n17), .C (x0), .Y (n122) );
  INVx1_ASAP7_75t_R    g0115( .A (n122), .Y (n123) );
  AND2x2_ASAP7_75t_R   g0116( .A (n121), .B (n123), .Y (y31) );
  NAND2x1_ASAP7_75t_R  g0117( .A (x0), .B (n17), .Y (n125) );
  AO21x1_ASAP7_75t_R   g0118( .A1 (n125), .A2 (n84), .B (n13), .Y (y32) );
  NOR2x1_ASAP7_75t_R   g0119( .A (x3), .B (x0), .Y (n127) );
  NOR2x1_ASAP7_75t_R   g0120( .A (x1), .B (x2), .Y (n128) );
  INVx1_ASAP7_75t_R    g0121( .A (n128), .Y (n129) );
  AND2x2_ASAP7_75t_R   g0122( .A (x3), .B (x0), .Y (n130) );
  AO21x1_ASAP7_75t_R   g0123( .A1 (x1), .A2 (x2), .B (n130), .Y (n131) );
  AO21x1_ASAP7_75t_R   g0124( .A1 (n127), .A2 (n129), .B (n131), .Y (y33) );
  AO21x1_ASAP7_75t_R   g0125( .A1 (n17), .A2 (x2), .B (n12), .Y (n133) );
  NAND2x1_ASAP7_75t_R  g0126( .A (n105), .B (n133), .Y (y34) );
  INVx1_ASAP7_75t_R    g0127( .A (n117), .Y (n135) );
  OA21x2_ASAP7_75t_R   g0128( .A1 (n103), .A2 (n116), .B (n135), .Y (y35) );
  NAND2x1_ASAP7_75t_R  g0129( .A (x2), .B (n17), .Y (n137) );
  AO21x1_ASAP7_75t_R   g0130( .A1 (n137), .A2 (x0), .B (n103), .Y (y36) );
  NOR2x1_ASAP7_75t_R   g0131( .A (x0), .B (x3), .Y (n139) );
  AND3x1_ASAP7_75t_R   g0132( .A (n139), .B (n15), .C (n16), .Y (n140) );
  NOR2x1_ASAP7_75t_R   g0133( .A (n12), .B (n111), .Y (n141) );
  OR3x1_ASAP7_75t_R    g0134( .A (n140), .B (n141), .C (n103), .Y (y37) );
  AND2x2_ASAP7_75t_R   g0135( .A (x0), .B (x1), .Y (n143) );
  INVx1_ASAP7_75t_R    g0136( .A (n143), .Y (n144) );
  AND2x2_ASAP7_75t_R   g0137( .A (x0), .B (x3), .Y (n145) );
  AO21x1_ASAP7_75t_R   g0138( .A1 (x1), .A2 (x2), .B (n145), .Y (n146) );
  AO21x1_ASAP7_75t_R   g0139( .A1 (n45), .A2 (n144), .B (n146), .Y (y38) );
  AO21x1_ASAP7_75t_R   g0140( .A1 (n15), .A2 (n16), .B (x3), .Y (n148) );
  AO21x1_ASAP7_75t_R   g0141( .A1 (n148), .A2 (x0), .B (n13), .Y (y39) );
  AO21x1_ASAP7_75t_R   g0142( .A1 (x2), .A2 (x1), .B (n130), .Y (y40) );
  AND3x1_ASAP7_75t_R   g0143( .A (n17), .B (x2), .C (x1), .Y (n151) );
  INVx1_ASAP7_75t_R    g0144( .A (n151), .Y (n152) );
  AO21x1_ASAP7_75t_R   g0145( .A1 (x1), .A2 (x2), .B (n17), .Y (n153) );
  AO21x1_ASAP7_75t_R   g0146( .A1 (n152), .A2 (n153), .B (x0), .Y (y41) );
  AO21x1_ASAP7_75t_R   g0147( .A1 (n15), .A2 (n16), .B (n12), .Y (n155) );
  INVx1_ASAP7_75t_R    g0148( .A (n155), .Y (y1081) );
  AND2x2_ASAP7_75t_R   g0149( .A (y25), .B (x3), .Y (n157) );
  NOR2x1_ASAP7_75t_R   g0150( .A (x3), .B (y25), .Y (n158) );
  OR3x1_ASAP7_75t_R    g0151( .A (y1081), .B (n157), .C (n158), .Y (y42) );
  NOR2x1_ASAP7_75t_R   g0152( .A (n51), .B (n85), .Y (n160) );
  OR3x1_ASAP7_75t_R    g0153( .A (n13), .B (n17), .C (x0), .Y (n161) );
  OA21x2_ASAP7_75t_R   g0154( .A1 (x3), .A2 (n160), .B (n161), .Y (y43) );
  INVx1_ASAP7_75t_R    g0155( .A (n137), .Y (n163) );
  INVx1_ASAP7_75t_R    g0156( .A (n72), .Y (n164) );
  OR3x1_ASAP7_75t_R    g0157( .A (n163), .B (n164), .C (n16), .Y (n165) );
  NAND2x1_ASAP7_75t_R  g0158( .A (n12), .B (n165), .Y (y44) );
  OR3x1_ASAP7_75t_R    g0159( .A (x0), .B (x3), .C (x2), .Y (n167) );
  AO21x1_ASAP7_75t_R   g0160( .A1 (n17), .A2 (n15), .B (n12), .Y (n168) );
  NAND2x1_ASAP7_75t_R  g0161( .A (n167), .B (n168), .Y (n169) );
  AO21x1_ASAP7_75t_R   g0162( .A1 (x1), .A2 (n9), .B (n169), .Y (y45) );
  AO21x1_ASAP7_75t_R   g0163( .A1 (x2), .A2 (x1), .B (n17), .Y (n171) );
  AO21x1_ASAP7_75t_R   g0164( .A1 (n148), .A2 (n171), .B (x0), .Y (y46) );
  INVx1_ASAP7_75t_R    g0165( .A (y863), .Y (n173) );
  AO21x1_ASAP7_75t_R   g0166( .A1 (n16), .A2 (n12), .B (n15), .Y (n174) );
  OR3x1_ASAP7_75t_R    g0167( .A (x1), .B (x0), .C (x2), .Y (n175) );
  AND3x1_ASAP7_75t_R   g0168( .A (n173), .B (n174), .C (n175), .Y (n176) );
  NAND2x1_ASAP7_75t_R  g0169( .A (x5), .B (n176), .Y (y47) );
  INVx1_ASAP7_75t_R    g0170( .A (n53), .Y (n178) );
  AO21x1_ASAP7_75t_R   g0171( .A1 (n178), .A2 (x0), .B (n65), .Y (y48) );
  AO21x1_ASAP7_75t_R   g0172( .A1 (n16), .A2 (x5), .B (n12), .Y (n180) );
  INVx1_ASAP7_75t_R    g0173( .A (n180), .Y (y772) );
  AND3x1_ASAP7_75t_R   g0174( .A (n51), .B (n12), .C (x5), .Y (n182) );
  OR3x1_ASAP7_75t_R    g0175( .A (n57), .B (y772), .C (n182), .Y (y49) );
  AND3x1_ASAP7_75t_R   g0176( .A (n16), .B (n12), .C (x3), .Y (n184) );
  AO21x1_ASAP7_75t_R   g0177( .A1 (x1), .A2 (x0), .B (x2), .Y (n185) );
  AND3x1_ASAP7_75t_R   g0178( .A (n16), .B (n12), .C (x2), .Y (n186) );
  INVx1_ASAP7_75t_R    g0179( .A (n186), .Y (n187) );
  OA21x2_ASAP7_75t_R   g0180( .A1 (n184), .A2 (n185), .B (n187), .Y (y50) );
  INVx1_ASAP7_75t_R    g0181( .A (n139), .Y (n189) );
  AND3x1_ASAP7_75t_R   g0182( .A (n129), .B (n189), .C (n113), .Y (y69) );
  AO21x1_ASAP7_75t_R   g0183( .A1 (x2), .A2 (x3), .B (x0), .Y (n191) );
  NOR2x1_ASAP7_75t_R   g0184( .A (x1), .B (n191), .Y (n192) );
  OR3x1_ASAP7_75t_R    g0185( .A (y69), .B (n45), .C (n192), .Y (y51) );
  OR3x1_ASAP7_75t_R    g0186( .A (n43), .B (n17), .C (n15), .Y (n194) );
  INVx1_ASAP7_75t_R    g0187( .A (n194), .Y (n195) );
  OR3x1_ASAP7_75t_R    g0188( .A (n195), .B (n143), .C (n192), .Y (y2991) );
  AO21x1_ASAP7_75t_R   g0189( .A1 (n15), .A2 (n17), .B (y2991), .Y (y52) );
  NAND2x1_ASAP7_75t_R  g0190( .A (n175), .B (n174), .Y (n198) );
  AO21x1_ASAP7_75t_R   g0191( .A1 (n174), .A2 (n175), .B (n17), .Y (n199) );
  OA21x2_ASAP7_75t_R   g0192( .A1 (n198), .A2 (x3), .B (n199), .Y (n200) );
  NAND2x1_ASAP7_75t_R  g0193( .A (n173), .B (n200), .Y (y53) );
  AO21x1_ASAP7_75t_R   g0194( .A1 (n12), .A2 (n17), .B (n15), .Y (n202) );
  INVx1_ASAP7_75t_R    g0195( .A (n202), .Y (n203) );
  AO21x1_ASAP7_75t_R   g0196( .A1 (x0), .A2 (x3), .B (x1), .Y (n204) );
  AO21x1_ASAP7_75t_R   g0197( .A1 (n12), .A2 (n15), .B (n17), .Y (n205) );
  AO21x1_ASAP7_75t_R   g0198( .A1 (x0), .A2 (x2), .B (x1), .Y (n206) );
  INVx1_ASAP7_75t_R    g0199( .A (n206), .Y (n207) );
  AO21x1_ASAP7_75t_R   g0200( .A1 (n205), .A2 (n207), .B (n143), .Y (n208) );
  AO21x1_ASAP7_75t_R   g0201( .A1 (n203), .A2 (n204), .B (n208), .Y (y54) );
  AO21x1_ASAP7_75t_R   g0202( .A1 (n15), .A2 (n17), .B (x1), .Y (n210) );
  AND2x2_ASAP7_75t_R   g0203( .A (x2), .B (x3), .Y (n211) );
  AO21x1_ASAP7_75t_R   g0204( .A1 (n210), .A2 (x0), .B (n211), .Y (n212) );
  AO21x1_ASAP7_75t_R   g0205( .A1 (n137), .A2 (n72), .B (x0), .Y (n213) );
  NOR2x1_ASAP7_75t_R   g0206( .A (x1), .B (n213), .Y (n214) );
  AO21x1_ASAP7_75t_R   g0207( .A1 (n46), .A2 (n212), .B (n214), .Y (y55) );
  AO21x1_ASAP7_75t_R   g0208( .A1 (x2), .A2 (x3), .B (y863), .Y (n216) );
  AND2x2_ASAP7_75t_R   g0209( .A (n137), .B (n72), .Y (n217) );
  INVx1_ASAP7_75t_R    g0210( .A (n217), .Y (n218) );
  NAND2x1_ASAP7_75t_R  g0211( .A (x1), .B (n12), .Y (n219) );
  AND2x2_ASAP7_75t_R   g0212( .A (n90), .B (n219), .Y (y435) );
  INVx1_ASAP7_75t_R    g0213( .A (y435), .Y (n221) );
  AND2x2_ASAP7_75t_R   g0214( .A (n218), .B (n221), .Y (n222) );
  AO21x1_ASAP7_75t_R   g0215( .A1 (n49), .A2 (n216), .B (n222), .Y (n223) );
  INVx1_ASAP7_75t_R    g0216( .A (n223), .Y (y56) );
  AND3x1_ASAP7_75t_R   g0217( .A (n173), .B (n174), .C (x5), .Y (n225) );
  INVx1_ASAP7_75t_R    g0218( .A (n225), .Y (y57) );
  NOR2x1_ASAP7_75t_R   g0219( .A (x1), .B (x0), .Y (n227) );
  INVx1_ASAP7_75t_R    g0220( .A (n227), .Y (n228) );
  AO21x1_ASAP7_75t_R   g0221( .A1 (y2079), .A2 (x2), .B (y863), .Y (y2770) );
  AO21x1_ASAP7_75t_R   g0222( .A1 (n97), .A2 (n228), .B (y2770), .Y (y58) );
  NOR2x1_ASAP7_75t_R   g0223( .A (x1), .B (x5), .Y (n231) );
  AO21x1_ASAP7_75t_R   g0224( .A1 (n231), .A2 (n12), .B (y863), .Y (n232) );
  OA21x2_ASAP7_75t_R   g0225( .A1 (x2), .A2 (n232), .B (n187), .Y (y59) );
  NAND2x1_ASAP7_75t_R  g0226( .A (n174), .B (n173), .Y (y60) );
  AND3x1_ASAP7_75t_R   g0227( .A (n17), .B (x1), .C (x2), .Y (n235) );
  INVx1_ASAP7_75t_R    g0228( .A (n235), .Y (n236) );
  AO21x1_ASAP7_75t_R   g0229( .A1 (n236), .A2 (n171), .B (y1081), .Y (y61) );
  NAND2x1_ASAP7_75t_R  g0230( .A (n128), .B (n125), .Y (n238) );
  AND2x2_ASAP7_75t_R   g0231( .A (y41), .B (n238), .Y (y62) );
  OA33x2_ASAP7_75t_R   g0232( .A1 (n16), .A2 (n137), .A3 (x0), .B1 (n139), .B2 (y1081), .B3 (n13), .Y (y63) );
  NOR2x1_ASAP7_75t_R   g0233( .A (x0), .B (x2), .Y (n241) );
  INVx1_ASAP7_75t_R    g0234( .A (n241), .Y (n242) );
  AND2x2_ASAP7_75t_R   g0235( .A (x1), .B (x3), .Y (n243) );
  NAND2x1_ASAP7_75t_R  g0236( .A (x2), .B (n12), .Y (n244) );
  AND2x2_ASAP7_75t_R   g0237( .A (n72), .B (n244), .Y (n245) );
  AO21x1_ASAP7_75t_R   g0238( .A1 (n242), .A2 (n243), .B (n245), .Y (y64) );
  AO21x1_ASAP7_75t_R   g0239( .A1 (n12), .A2 (x3), .B (n15), .Y (n247) );
  AND2x2_ASAP7_75t_R   g0240( .A (n247), .B (x1), .Y (n248) );
  OR3x1_ASAP7_75t_R    g0241( .A (n143), .B (n17), .C (x2), .Y (n249) );
  OA21x2_ASAP7_75t_R   g0242( .A1 (x0), .A2 (n248), .B (n249), .Y (y65) );
  AO21x1_ASAP7_75t_R   g0243( .A1 (n17), .A2 (n241), .B (y69), .Y (y66) );
  AO21x1_ASAP7_75t_R   g0244( .A1 (n16), .A2 (n17), .B (x2), .Y (n252) );
  AO21x1_ASAP7_75t_R   g0245( .A1 (x1), .A2 (x3), .B (n15), .Y (n253) );
  AO21x1_ASAP7_75t_R   g0246( .A1 (n252), .A2 (n253), .B (y1081), .Y (y67) );
  OR3x1_ASAP7_75t_R    g0247( .A (x0), .B (x1), .C (x3), .Y (n255) );
  INVx1_ASAP7_75t_R    g0248( .A (n255), .Y (n256) );
  AO21x1_ASAP7_75t_R   g0249( .A1 (n15), .A2 (n256), .B (y69), .Y (y68) );
  AO21x1_ASAP7_75t_R   g0250( .A1 (n16), .A2 (n12), .B (n17), .Y (n258) );
  INVx1_ASAP7_75t_R    g0251( .A (n258), .Y (n259) );
  AO21x1_ASAP7_75t_R   g0252( .A1 (x1), .A2 (x0), .B (x3), .Y (n260) );
  INVx1_ASAP7_75t_R    g0253( .A (n260), .Y (n261) );
  AND3x1_ASAP7_75t_R   g0254( .A (x1), .B (x0), .C (x2), .Y (n262) );
  AO21x1_ASAP7_75t_R   g0255( .A1 (n174), .A2 (n261), .B (n262), .Y (n263) );
  AO21x1_ASAP7_75t_R   g0256( .A1 (n259), .A2 (n185), .B (n263), .Y (y70) );
  AO21x1_ASAP7_75t_R   g0257( .A1 (n128), .A2 (n17), .B (n143), .Y (n265) );
  AO21x1_ASAP7_75t_R   g0258( .A1 (n76), .A2 (y9), .B (n265), .Y (y71) );
  AO21x1_ASAP7_75t_R   g0259( .A1 (n17), .A2 (n15), .B (x1), .Y (n267) );
  AND2x2_ASAP7_75t_R   g0260( .A (n267), .B (x0), .Y (n268) );
  AO21x1_ASAP7_75t_R   g0261( .A1 (y9), .A2 (n76), .B (n268), .Y (y72) );
  AO21x1_ASAP7_75t_R   g0262( .A1 (y9), .A2 (n76), .B (n143), .Y (y73) );
  INVx1_ASAP7_75t_R    g0263( .A (n185), .Y (n271) );
  AO21x1_ASAP7_75t_R   g0264( .A1 (x0), .A2 (n103), .B (n271), .Y (n272) );
  OR3x1_ASAP7_75t_R    g0265( .A (y863), .B (n17), .C (x2), .Y (n273) );
  OA21x2_ASAP7_75t_R   g0266( .A1 (n259), .A2 (n272), .B (n273), .Y (y74) );
  INVx1_ASAP7_75t_R    g0267( .A (n205), .Y (n275) );
  AND2x2_ASAP7_75t_R   g0268( .A (x0), .B (x2), .Y (n276) );
  AO21x1_ASAP7_75t_R   g0269( .A1 (x1), .A2 (n276), .B (n128), .Y (n277) );
  AND2x2_ASAP7_75t_R   g0270( .A (n277), .B (n17), .Y (n278) );
  AO21x1_ASAP7_75t_R   g0271( .A1 (n206), .A2 (n275), .B (n278), .Y (y75) );
  NAND2x1_ASAP7_75t_R  g0272( .A (n19), .B (n18), .Y (n280) );
  AO32x1_ASAP7_75t_R   g0273( .A1 (x2), .A2 (x1), .A3 (n189), .B1 (x0), .B2 (n280), .Y (y76) );
  AO21x1_ASAP7_75t_R   g0274( .A1 (n17), .A2 (n15), .B (n43), .Y (n282) );
  AO21x1_ASAP7_75t_R   g0275( .A1 (n144), .A2 (n77), .B (n282), .Y (n283) );
  INVx1_ASAP7_75t_R    g0276( .A (n283), .Y (y77) );
  AO21x1_ASAP7_75t_R   g0277( .A1 (n22), .A2 (n17), .B (x5), .Y (n285) );
  INVx1_ASAP7_75t_R    g0278( .A (n285), .Y (n286) );
  AO21x1_ASAP7_75t_R   g0279( .A1 (x4), .A2 (x3), .B (y2079), .Y (n287) );
  INVx1_ASAP7_75t_R    g0280( .A (n287), .Y (n288) );
  OR3x1_ASAP7_75t_R    g0281( .A (n286), .B (n288), .C (x0), .Y (y78) );
  NAND2x1_ASAP7_75t_R  g0282( .A (x4), .B (n17), .Y (n290) );
  INVx1_ASAP7_75t_R    g0283( .A (n290), .Y (n291) );
  AO21x1_ASAP7_75t_R   g0284( .A1 (x4), .A2 (x5), .B (n17), .Y (n292) );
  INVx1_ASAP7_75t_R    g0285( .A (n292), .Y (n293) );
  OR3x1_ASAP7_75t_R    g0286( .A (n291), .B (n293), .C (n58), .Y (y79) );
  AO21x1_ASAP7_75t_R   g0287( .A1 (x5), .A2 (x4), .B (n17), .Y (n295) );
  INVx1_ASAP7_75t_R    g0288( .A (n295), .Y (n296) );
  AND3x1_ASAP7_75t_R   g0289( .A (n17), .B (x5), .C (x4), .Y (n297) );
  OR3x1_ASAP7_75t_R    g0290( .A (n296), .B (n297), .C (x0), .Y (y80) );
  NAND2x1_ASAP7_75t_R  g0291( .A (x4), .B (n12), .Y (n299) );
  AND3x1_ASAP7_75t_R   g0292( .A (n22), .B (x5), .C (x0), .Y (n300) );
  INVx1_ASAP7_75t_R    g0293( .A (n300), .Y (n301) );
  NAND2x1_ASAP7_75t_R  g0294( .A (x5), .B (n12), .Y (y3852) );
  AND3x1_ASAP7_75t_R   g0295( .A (n12), .B (n17), .C (x5), .Y (n303) );
  AO21x1_ASAP7_75t_R   g0296( .A1 (y3852), .A2 (x3), .B (n303), .Y (n304) );
  AO21x1_ASAP7_75t_R   g0297( .A1 (n299), .A2 (n301), .B (n304), .Y (y81) );
  AND3x1_ASAP7_75t_R   g0298( .A (n12), .B (n22), .C (x5), .Y (n306) );
  AO21x1_ASAP7_75t_R   g0299( .A1 (n22), .A2 (x5), .B (n12), .Y (n307) );
  INVx1_ASAP7_75t_R    g0300( .A (n307), .Y (n308) );
  OR3x1_ASAP7_75t_R    g0301( .A (n304), .B (n306), .C (n308), .Y (y82) );
  NAND2x1_ASAP7_75t_R  g0302( .A (x0), .B (n22), .Y (n310) );
  AO21x1_ASAP7_75t_R   g0303( .A1 (n299), .A2 (n310), .B (n304), .Y (y83) );
  NAND2x1_ASAP7_75t_R  g0304( .A (x1), .B (y2079), .Y (n312) );
  NOR2x1_ASAP7_75t_R   g0305( .A (n310), .B (n312), .Y (y3428) );
  NOR2x1_ASAP7_75t_R   g0306( .A (n26), .B (y3428), .Y (y84) );
  NOR2x1_ASAP7_75t_R   g0307( .A (x0), .B (x4), .Y (n315) );
  NAND2x1_ASAP7_75t_R  g0308( .A (x3), .B (y2079), .Y (n316) );
  NAND2x1_ASAP7_75t_R  g0309( .A (n315), .B (n316), .Y (n317) );
  INVx1_ASAP7_75t_R    g0310( .A (n317), .Y (n318) );
  NAND2x1_ASAP7_75t_R  g0311( .A (x5), .B (n17), .Y (n319) );
  AO21x1_ASAP7_75t_R   g0312( .A1 (n316), .A2 (n319), .B (n22), .Y (n320) );
  INVx1_ASAP7_75t_R    g0313( .A (n320), .Y (n321) );
  AO21x1_ASAP7_75t_R   g0314( .A1 (n17), .A2 (x5), .B (n12), .Y (n322) );
  INVx1_ASAP7_75t_R    g0315( .A (n322), .Y (n323) );
  OR3x1_ASAP7_75t_R    g0316( .A (n318), .B (n321), .C (n323), .Y (y85) );
  AND2x2_ASAP7_75t_R   g0317( .A (x4), .B (x3), .Y (n325) );
  OR3x1_ASAP7_75t_R    g0318( .A (n325), .B (y2079), .C (x0), .Y (n326) );
  INVx1_ASAP7_75t_R    g0319( .A (n326), .Y (n327) );
  AO21x1_ASAP7_75t_R   g0320( .A1 (n22), .A2 (n17), .B (n12), .Y (n328) );
  INVx1_ASAP7_75t_R    g0321( .A (n328), .Y (n329) );
  AO21x1_ASAP7_75t_R   g0322( .A1 (x4), .A2 (x3), .B (x0), .Y (n330) );
  NAND2x1_ASAP7_75t_R  g0323( .A (y2079), .B (n330), .Y (n331) );
  INVx1_ASAP7_75t_R    g0324( .A (n331), .Y (n332) );
  OR3x1_ASAP7_75t_R    g0325( .A (n327), .B (n329), .C (n332), .Y (y86) );
  AO21x1_ASAP7_75t_R   g0326( .A1 (x3), .A2 (x4), .B (n12), .Y (n334) );
  AND3x1_ASAP7_75t_R   g0327( .A (x5), .B (x3), .C (x4), .Y (n335) );
  INVx1_ASAP7_75t_R    g0328( .A (n335), .Y (n336) );
  NOR2x1_ASAP7_75t_R   g0329( .A (x3), .B (x4), .Y (n337) );
  OR3x1_ASAP7_75t_R    g0330( .A (n337), .B (y2079), .C (n12), .Y (n338) );
  INVx1_ASAP7_75t_R    g0331( .A (n338), .Y (n339) );
  AO21x1_ASAP7_75t_R   g0332( .A1 (n334), .A2 (n336), .B (n339), .Y (y87) );
  AO21x1_ASAP7_75t_R   g0333( .A1 (n12), .A2 (y2079), .B (n22), .Y (n341) );
  INVx1_ASAP7_75t_R    g0334( .A (n341), .Y (n342) );
  OR3x1_ASAP7_75t_R    g0335( .A (x0), .B (x4), .C (x5), .Y (n343) );
  INVx1_ASAP7_75t_R    g0336( .A (n343), .Y (n344) );
  OA33x2_ASAP7_75t_R   g0337( .A1 (x3), .A2 (n342), .A3 (n344), .B1 (n17), .B2 (n22), .B3 (y3852), .Y (y88) );
  NAND2x1_ASAP7_75t_R  g0338( .A (n12), .B (n287), .Y (n346) );
  NOR2x1_ASAP7_75t_R   g0339( .A (x4), .B (x3), .Y (n347) );
  INVx1_ASAP7_75t_R    g0340( .A (n347), .Y (n348) );
  AND3x1_ASAP7_75t_R   g0341( .A (y2079), .B (x3), .C (x4), .Y (n349) );
  AO21x1_ASAP7_75t_R   g0342( .A1 (n346), .A2 (n348), .B (n349), .Y (y89) );
  AO21x1_ASAP7_75t_R   g0343( .A1 (y2079), .A2 (x0), .B (x3), .Y (n351) );
  NAND2x1_ASAP7_75t_R  g0344( .A (x0), .B (y2079), .Y (n352) );
  AO21x1_ASAP7_75t_R   g0345( .A1 (n12), .A2 (x5), .B (n17), .Y (n353) );
  INVx1_ASAP7_75t_R    g0346( .A (n353), .Y (n354) );
  AO221x2_ASAP7_75t_R  g0347( .A1 (n22), .A2 (n351), .B1 (n352), .B2 (n291), .C (n354), .Y (y90) );
  AO21x1_ASAP7_75t_R   g0348( .A1 (n12), .A2 (n17), .B (x5), .Y (n356) );
  NAND2x1_ASAP7_75t_R  g0349( .A (x4), .B (n356), .Y (n357) );
  INVx1_ASAP7_75t_R    g0350( .A (n357), .Y (n358) );
  AO21x1_ASAP7_75t_R   g0351( .A1 (n358), .A2 (n84), .B (n293), .Y (y91) );
  NAND2x1_ASAP7_75t_R  g0352( .A (x3), .B (n22), .Y (n360) );
  AO21x1_ASAP7_75t_R   g0353( .A1 (n290), .A2 (n360), .B (y2079), .Y (n361) );
  INVx1_ASAP7_75t_R    g0354( .A (n361), .Y (n362) );
  NOR2x1_ASAP7_75t_R   g0355( .A (x0), .B (x5), .Y (n363) );
  AND2x2_ASAP7_75t_R   g0356( .A (n360), .B (n363), .Y (n364) );
  OR3x1_ASAP7_75t_R    g0357( .A (n362), .B (n364), .C (n145), .Y (y92) );
  AO21x1_ASAP7_75t_R   g0358( .A1 (n22), .A2 (x3), .B (y2079), .Y (n366) );
  AO21x1_ASAP7_75t_R   g0359( .A1 (x4), .A2 (n17), .B (n366), .Y (n367) );
  AND2x2_ASAP7_75t_R   g0360( .A (x3), .B (x5), .Y (n368) );
  INVx1_ASAP7_75t_R    g0361( .A (n368), .Y (n369) );
  AO21x1_ASAP7_75t_R   g0362( .A1 (n17), .A2 (y2079), .B (n22), .Y (n370) );
  AO21x1_ASAP7_75t_R   g0363( .A1 (n369), .A2 (n370), .B (n12), .Y (n371) );
  INVx1_ASAP7_75t_R    g0364( .A (n371), .Y (n372) );
  AO21x1_ASAP7_75t_R   g0365( .A1 (n328), .A2 (n367), .B (n372), .Y (y93) );
  AND3x1_ASAP7_75t_R   g0366( .A (n12), .B (x4), .C (x3), .Y (n374) );
  NOR2x1_ASAP7_75t_R   g0367( .A (n347), .B (n374), .Y (n375) );
  NOR2x1_ASAP7_75t_R   g0368( .A (x5), .B (n139), .Y (n376) );
  AND2x2_ASAP7_75t_R   g0369( .A (n360), .B (n290), .Y (n377) );
  INVx1_ASAP7_75t_R    g0370( .A (n377), .Y (n378) );
  AND3x1_ASAP7_75t_R   g0371( .A (n378), .B (y2079), .C (x0), .Y (y2376) );
  INVx1_ASAP7_75t_R    g0372( .A (y2376), .Y (n380) );
  OA21x2_ASAP7_75t_R   g0373( .A1 (n375), .A2 (n376), .B (n380), .Y (y94) );
  INVx1_ASAP7_75t_R    g0374( .A (n325), .Y (n382) );
  AND3x1_ASAP7_75t_R   g0375( .A (x0), .B (x4), .C (x3), .Y (n383) );
  AO21x1_ASAP7_75t_R   g0376( .A1 (n382), .A2 (x5), .B (n383), .Y (n384) );
  AO21x1_ASAP7_75t_R   g0377( .A1 (n384), .A2 (n348), .B (n363), .Y (y95) );
  AND3x1_ASAP7_75t_R   g0378( .A (n12), .B (x4), .C (x5), .Y (n386) );
  INVx1_ASAP7_75t_R    g0379( .A (n386), .Y (n387) );
  NAND2x1_ASAP7_75t_R  g0380( .A (x4), .B (y2079), .Y (n388) );
  AND3x1_ASAP7_75t_R   g0381( .A (n388), .B (n28), .C (n17), .Y (n389) );
  AO21x1_ASAP7_75t_R   g0382( .A1 (n387), .A2 (x3), .B (n389), .Y (y96) );
  AO21x1_ASAP7_75t_R   g0383( .A1 (y2079), .A2 (n22), .B (x3), .Y (n391) );
  AND2x2_ASAP7_75t_R   g0384( .A (x5), .B (x4), .Y (n392) );
  INVx1_ASAP7_75t_R    g0385( .A (n392), .Y (y3293) );
  AO21x1_ASAP7_75t_R   g0386( .A1 (y3293), .A2 (x3), .B (n297), .Y (y2578) );
  AO21x1_ASAP7_75t_R   g0387( .A1 (x0), .A2 (n391), .B (y2578), .Y (y97) );
  AND2x2_ASAP7_75t_R   g0388( .A (n388), .B (n28), .Y (n396) );
  AO21x1_ASAP7_75t_R   g0389( .A1 (n17), .A2 (x5), .B (x0), .Y (n397) );
  AO21x1_ASAP7_75t_R   g0390( .A1 (n388), .A2 (n28), .B (n17), .Y (n398) );
  INVx1_ASAP7_75t_R    g0391( .A (n398), .Y (n399) );
  AO21x1_ASAP7_75t_R   g0392( .A1 (n396), .A2 (n397), .B (n399), .Y (y98) );
  INVx1_ASAP7_75t_R    g0393( .A (n337), .Y (n401) );
  OR3x1_ASAP7_75t_R    g0394( .A (n17), .B (n22), .C (x0), .Y (n402) );
  AND2x2_ASAP7_75t_R   g0395( .A (x3), .B (x4), .Y (n403) );
  AO21x1_ASAP7_75t_R   g0396( .A1 (n12), .A2 (n22), .B (n403), .Y (n404) );
  AO32x1_ASAP7_75t_R   g0397( .A1 (x5), .A2 (n401), .A3 (n402), .B1 (y2079), .B2 (n404), .Y (y99) );
  AO21x1_ASAP7_75t_R   g0398( .A1 (n17), .A2 (n22), .B (y2079), .Y (n406) );
  INVx1_ASAP7_75t_R    g0399( .A (n406), .Y (n407) );
  AO21x1_ASAP7_75t_R   g0400( .A1 (n22), .A2 (x0), .B (n17), .Y (n408) );
  INVx1_ASAP7_75t_R    g0401( .A (n408), .Y (n409) );
  AND3x1_ASAP7_75t_R   g0402( .A (n12), .B (x5), .C (x4), .Y (n410) );
  NAND2x1_ASAP7_75t_R  g0403( .A (x3), .B (n410), .Y (n411) );
  OA21x2_ASAP7_75t_R   g0404( .A1 (n407), .A2 (n409), .B (n411), .Y (y100) );
  INVx1_ASAP7_75t_R    g0405( .A (n374), .Y (n413) );
  AO21x1_ASAP7_75t_R   g0406( .A1 (n413), .A2 (n348), .B (y2079), .Y (y3134) );
  AO21x1_ASAP7_75t_R   g0407( .A1 (n17), .A2 (x0), .B (x4), .Y (n415) );
  AO21x1_ASAP7_75t_R   g0408( .A1 (n290), .A2 (n415), .B (x5), .Y (n416) );
  AND2x2_ASAP7_75t_R   g0409( .A (y3134), .B (n416), .Y (y101) );
  NOR2x1_ASAP7_75t_R   g0410( .A (x5), .B (x4), .Y (n418) );
  INVx1_ASAP7_75t_R    g0411( .A (n418), .Y (n419) );
  INVx1_ASAP7_75t_R    g0412( .A (n410), .Y (y103) );
  INVx1_ASAP7_75t_R    g0413( .A (n319), .Y (n421) );
  AO32x1_ASAP7_75t_R   g0414( .A1 (n419), .A2 (y103), .A3 (x3), .B1 (n421), .B2 (x4), .Y (y102) );
  AO21x1_ASAP7_75t_R   g0415( .A1 (x4), .A2 (y2079), .B (n23), .Y (y104) );
  INVx1_ASAP7_75t_R    g0416( .A (n396), .Y (y3758) );
  AND3x1_ASAP7_75t_R   g0417( .A (n12), .B (y2079), .C (x3), .Y (n425) );
  AO21x1_ASAP7_75t_R   g0418( .A1 (y2079), .A2 (x3), .B (n12), .Y (n426) );
  INVx1_ASAP7_75t_R    g0419( .A (n426), .Y (n427) );
  OR3x1_ASAP7_75t_R    g0420( .A (y3758), .B (n425), .C (n427), .Y (y105) );
  AO21x1_ASAP7_75t_R   g0421( .A1 (x5), .A2 (x4), .B (x0), .Y (n429) );
  AO21x1_ASAP7_75t_R   g0422( .A1 (y2079), .A2 (n22), .B (n12), .Y (n430) );
  NAND2x1_ASAP7_75t_R  g0423( .A (n429), .B (n430), .Y (y106) );
  OR3x1_ASAP7_75t_R    g0424( .A (n139), .B (x4), .C (x5), .Y (n432) );
  AND2x2_ASAP7_75t_R   g0425( .A (y103), .B (n432), .Y (y107) );
  AO21x1_ASAP7_75t_R   g0426( .A1 (y2079), .A2 (n22), .B (n410), .Y (n434) );
  INVx1_ASAP7_75t_R    g0427( .A (n434), .Y (y108) );
  NAND2x1_ASAP7_75t_R  g0428( .A (x1), .B (n22), .Y (n436) );
  INVx1_ASAP7_75t_R    g0429( .A (n436), .Y (n437) );
  OR3x1_ASAP7_75t_R    g0430( .A (n437), .B (y2079), .C (x0), .Y (y109) );
  AO21x1_ASAP7_75t_R   g0431( .A1 (n22), .A2 (y2079), .B (n12), .Y (n439) );
  INVx1_ASAP7_75t_R    g0432( .A (n439), .Y (n440) );
  OR3x1_ASAP7_75t_R    g0433( .A (n437), .B (n440), .C (n363), .Y (y110) );
  AND3x1_ASAP7_75t_R   g0434( .A (n22), .B (x5), .C (x1), .Y (n442) );
  AO21x1_ASAP7_75t_R   g0435( .A1 (n436), .A2 (y2079), .B (x0), .Y (n443) );
  AND3x1_ASAP7_75t_R   g0436( .A (y2466), .B (n16), .C (x0), .Y (n444) );
  INVx1_ASAP7_75t_R    g0437( .A (n444), .Y (n445) );
  OA21x2_ASAP7_75t_R   g0438( .A1 (n442), .A2 (n443), .B (n445), .Y (y111) );
  AO21x1_ASAP7_75t_R   g0439( .A1 (n12), .A2 (x5), .B (y2466), .Y (n447) );
  OR3x1_ASAP7_75t_R    g0440( .A (n363), .B (n16), .C (x4), .Y (n448) );
  NAND2x1_ASAP7_75t_R  g0441( .A (n447), .B (n448), .Y (y112) );
  AND3x1_ASAP7_75t_R   g0442( .A (n22), .B (y2079), .C (x0), .Y (n450) );
  INVx1_ASAP7_75t_R    g0443( .A (n450), .Y (n451) );
  AND2x2_ASAP7_75t_R   g0444( .A (y109), .B (n451), .Y (y113) );
  OR3x1_ASAP7_75t_R    g0445( .A (n43), .B (x5), .C (x4), .Y (n453) );
  AND2x2_ASAP7_75t_R   g0446( .A (y109), .B (n453), .Y (y114) );
  INVx1_ASAP7_75t_R    g0447( .A (y2466), .Y (n455) );
  AND2x2_ASAP7_75t_R   g0448( .A (y109), .B (n455), .Y (y115) );
  AO21x1_ASAP7_75t_R   g0449( .A1 (y2079), .A2 (n22), .B (x1), .Y (n457) );
  AO21x1_ASAP7_75t_R   g0450( .A1 (y3293), .A2 (n457), .B (x0), .Y (y116) );
  AO21x1_ASAP7_75t_R   g0451( .A1 (x5), .A2 (x4), .B (n16), .Y (n459) );
  NAND2x1_ASAP7_75t_R  g0452( .A (n12), .B (n459), .Y (y117) );
  NAND2x1_ASAP7_75t_R  g0453( .A (n459), .B (n430), .Y (y118) );
  AND3x1_ASAP7_75t_R   g0454( .A (n22), .B (y2079), .C (x1), .Y (n462) );
  AO21x1_ASAP7_75t_R   g0455( .A1 (n22), .A2 (x1), .B (y2079), .Y (n463) );
  INVx1_ASAP7_75t_R    g0456( .A (n463), .Y (n464) );
  NOR2x1_ASAP7_75t_R   g0457( .A (n462), .B (n464), .Y (n465) );
  NAND2x1_ASAP7_75t_R  g0458( .A (x4), .B (n16), .Y (n466) );
  AO21x1_ASAP7_75t_R   g0459( .A1 (n465), .A2 (n466), .B (x0), .Y (y119) );
  AND3x1_ASAP7_75t_R   g0460( .A (y2079), .B (n22), .C (x1), .Y (n468) );
  INVx1_ASAP7_75t_R    g0461( .A (n468), .Y (n469) );
  AND2x2_ASAP7_75t_R   g0462( .A (y116), .B (n469), .Y (y120) );
  OR3x1_ASAP7_75t_R    g0463( .A (n43), .B (x4), .C (x5), .Y (n471) );
  AND2x2_ASAP7_75t_R   g0464( .A (y116), .B (n471), .Y (y121) );
  AO21x1_ASAP7_75t_R   g0465( .A1 (n12), .A2 (y2079), .B (x4), .Y (n473) );
  INVx1_ASAP7_75t_R    g0466( .A (n473), .Y (n474) );
  OR3x1_ASAP7_75t_R    g0467( .A (x1), .B (x4), .C (x5), .Y (n475) );
  INVx1_ASAP7_75t_R    g0468( .A (n475), .Y (n476) );
  AO221x2_ASAP7_75t_R  g0469( .A1 (x4), .A2 (y3852), .B1 (n90), .B2 (n474), .C (n476), .Y (y122) );
  AND3x1_ASAP7_75t_R   g0470( .A (n16), .B (n22), .C (x5), .Y (n478) );
  NOR2x1_ASAP7_75t_R   g0471( .A (n12), .B (n478), .Y (n479) );
  AO21x1_ASAP7_75t_R   g0472( .A1 (y3758), .A2 (n12), .B (n479), .Y (y123) );
  INVx1_ASAP7_75t_R    g0473( .A (y3852), .Y (n481) );
  AO21x1_ASAP7_75t_R   g0474( .A1 (x0), .A2 (x1), .B (x4), .Y (n482) );
  OA21x2_ASAP7_75t_R   g0475( .A1 (n481), .A2 (n482), .B (n387), .Y (y124) );
  AO21x1_ASAP7_75t_R   g0476( .A1 (x0), .A2 (x1), .B (x5), .Y (n484) );
  INVx1_ASAP7_75t_R    g0477( .A (n484), .Y (n485) );
  AO21x1_ASAP7_75t_R   g0478( .A1 (x1), .A2 (n58), .B (n485), .Y (n486) );
  AO21x1_ASAP7_75t_R   g0479( .A1 (n299), .A2 (n310), .B (n486), .Y (y125) );
  AO21x1_ASAP7_75t_R   g0480( .A1 (n12), .A2 (x5), .B (x1), .Y (n488) );
  AO21x1_ASAP7_75t_R   g0481( .A1 (x0), .A2 (x4), .B (y2079), .Y (n489) );
  AO21x1_ASAP7_75t_R   g0482( .A1 (n16), .A2 (x0), .B (x4), .Y (n490) );
  AO32x1_ASAP7_75t_R   g0483( .A1 (n488), .A2 (n352), .A3 (n22), .B1 (n489), .B2 (n490), .Y (y126) );
  AO21x1_ASAP7_75t_R   g0484( .A1 (n12), .A2 (x5), .B (n22), .Y (n492) );
  INVx1_ASAP7_75t_R    g0485( .A (n492), .Y (n493) );
  AO21x1_ASAP7_75t_R   g0486( .A1 (n29), .A2 (n90), .B (n493), .Y (y127) );
  INVx1_ASAP7_75t_R    g0487( .A (n312), .Y (n495) );
  OR3x1_ASAP7_75t_R    g0488( .A (n495), .B (n22), .C (x0), .Y (n496) );
  NAND2x1_ASAP7_75t_R  g0489( .A (x5), .B (n16), .Y (n497) );
  AO21x1_ASAP7_75t_R   g0490( .A1 (n312), .A2 (n497), .B (n310), .Y (n498) );
  AND2x2_ASAP7_75t_R   g0491( .A (n496), .B (n498), .Y (y128) );
  AO21x1_ASAP7_75t_R   g0492( .A1 (y2079), .A2 (x1), .B (x0), .Y (y195) );
  AO21x1_ASAP7_75t_R   g0493( .A1 (n16), .A2 (y2079), .B (x4), .Y (n501) );
  AO21x1_ASAP7_75t_R   g0494( .A1 (x0), .A2 (n16), .B (n28), .Y (n502) );
  INVx1_ASAP7_75t_R    g0495( .A (n502), .Y (n503) );
  AO21x1_ASAP7_75t_R   g0496( .A1 (y195), .A2 (n501), .B (n503), .Y (y129) );
  OR3x1_ASAP7_75t_R    g0497( .A (n392), .B (n12), .C (x1), .Y (n505) );
  AND2x2_ASAP7_75t_R   g0498( .A (y103), .B (n505), .Y (y130) );
  AO21x1_ASAP7_75t_R   g0499( .A1 (n12), .A2 (x4), .B (x1), .Y (n507) );
  AO21x1_ASAP7_75t_R   g0500( .A1 (n310), .A2 (x5), .B (n507), .Y (n508) );
  AND2x2_ASAP7_75t_R   g0501( .A (n508), .B (n387), .Y (y131) );
  AO21x1_ASAP7_75t_R   g0502( .A1 (n12), .A2 (n22), .B (y2079), .Y (n510) );
  AO21x1_ASAP7_75t_R   g0503( .A1 (x0), .A2 (x4), .B (x1), .Y (n511) );
  INVx1_ASAP7_75t_R    g0504( .A (n511), .Y (n512) );
  AO21x1_ASAP7_75t_R   g0505( .A1 (x4), .A2 (x5), .B (x1), .Y (n513) );
  AND2x2_ASAP7_75t_R   g0506( .A (y104), .B (n513), .Y (y698) );
  AO21x1_ASAP7_75t_R   g0507( .A1 (n510), .A2 (n512), .B (y698), .Y (y132) );
  AO21x1_ASAP7_75t_R   g0508( .A1 (n469), .A2 (y3293), .B (x0), .Y (n516) );
  AND2x2_ASAP7_75t_R   g0509( .A (n516), .B (n505), .Y (y133) );
  AND2x2_ASAP7_75t_R   g0510( .A (x4), .B (x5), .Y (n518) );
  OR3x1_ASAP7_75t_R    g0511( .A (n518), .B (n12), .C (x1), .Y (n519) );
  AND2x2_ASAP7_75t_R   g0512( .A (y104), .B (n519), .Y (y134) );
  AO21x1_ASAP7_75t_R   g0513( .A1 (x5), .A2 (x4), .B (n143), .Y (n521) );
  INVx1_ASAP7_75t_R    g0514( .A (n521), .Y (n522) );
  AO21x1_ASAP7_75t_R   g0515( .A1 (y2079), .A2 (n22), .B (n16), .Y (n523) );
  AO21x1_ASAP7_75t_R   g0516( .A1 (y3293), .A2 (n523), .B (n12), .Y (n524) );
  INVx1_ASAP7_75t_R    g0517( .A (n524), .Y (n525) );
  AO21x1_ASAP7_75t_R   g0518( .A1 (n430), .A2 (n522), .B (n525), .Y (y135) );
  NOR2x1_ASAP7_75t_R   g0519( .A (x1), .B (x4), .Y (n527) );
  NOR2x1_ASAP7_75t_R   g0520( .A (n527), .B (n386), .Y (y136) );
  INVx1_ASAP7_75t_R    g0521( .A (n388), .Y (n529) );
  NOR2x1_ASAP7_75t_R   g0522( .A (n12), .B (n231), .Y (n530) );
  OR3x1_ASAP7_75t_R    g0523( .A (n529), .B (n29), .C (n530), .Y (y137) );
  AND3x1_ASAP7_75t_R   g0524( .A (n315), .B (y2079), .C (x1), .Y (n532) );
  INVx1_ASAP7_75t_R    g0525( .A (n532), .Y (n533) );
  INVx1_ASAP7_75t_R    g0526( .A (n527), .Y (n534) );
  AO21x1_ASAP7_75t_R   g0527( .A1 (n534), .A2 (n299), .B (y2079), .Y (y250) );
  AND2x2_ASAP7_75t_R   g0528( .A (n533), .B (y250), .Y (y138) );
  AND2x2_ASAP7_75t_R   g0529( .A (x0), .B (x4), .Y (n537) );
  AO21x1_ASAP7_75t_R   g0530( .A1 (n12), .A2 (y2079), .B (n537), .Y (n538) );
  INVx1_ASAP7_75t_R    g0531( .A (n448), .Y (n539) );
  AO21x1_ASAP7_75t_R   g0532( .A1 (n436), .A2 (n538), .B (n539), .Y (y139) );
  AO21x1_ASAP7_75t_R   g0533( .A1 (n12), .A2 (y2079), .B (n16), .Y (n541) );
  INVx1_ASAP7_75t_R    g0534( .A (n541), .Y (n542) );
  OA21x2_ASAP7_75t_R   g0535( .A1 (x4), .A2 (n542), .B (n387), .Y (y140) );
  AND2x2_ASAP7_75t_R   g0536( .A (x1), .B (x5), .Y (n544) );
  AO21x1_ASAP7_75t_R   g0537( .A1 (n544), .A2 (n22), .B (n538), .Y (y141) );
  INVx1_ASAP7_75t_R    g0538( .A (n462), .Y (n546) );
  AND2x2_ASAP7_75t_R   g0539( .A (y250), .B (n546), .Y (y142) );
  AO21x1_ASAP7_75t_R   g0540( .A1 (n489), .A2 (n490), .B (n442), .Y (y143) );
  AND2x2_ASAP7_75t_R   g0541( .A (n436), .B (n363), .Y (n549) );
  OR3x1_ASAP7_75t_R    g0542( .A (n549), .B (n442), .C (n537), .Y (y144) );
  AO21x1_ASAP7_75t_R   g0543( .A1 (x1), .A2 (x5), .B (x4), .Y (n551) );
  INVx1_ASAP7_75t_R    g0544( .A (n551), .Y (n552) );
  NOR2x1_ASAP7_75t_R   g0545( .A (n552), .B (n386), .Y (y145) );
  AO21x1_ASAP7_75t_R   g0546( .A1 (x4), .A2 (x5), .B (n16), .Y (n554) );
  NAND2x1_ASAP7_75t_R  g0547( .A (n554), .B (n307), .Y (y146) );
  INVx1_ASAP7_75t_R    g0548( .A (n518), .Y (n556) );
  AO21x1_ASAP7_75t_R   g0549( .A1 (n556), .A2 (x1), .B (n537), .Y (y147) );
  AO21x1_ASAP7_75t_R   g0550( .A1 (n12), .A2 (x1), .B (x5), .Y (n558) );
  INVx1_ASAP7_75t_R    g0551( .A (n558), .Y (n559) );
  OA21x2_ASAP7_75t_R   g0552( .A1 (n559), .A2 (n551), .B (n496), .Y (y148) );
  AO21x1_ASAP7_75t_R   g0553( .A1 (n388), .A2 (n28), .B (n16), .Y (n561) );
  NAND2x1_ASAP7_75t_R  g0554( .A (n307), .B (n561), .Y (y149) );
  AND3x1_ASAP7_75t_R   g0555( .A (n12), .B (y2079), .C (x1), .Y (n563) );
  INVx1_ASAP7_75t_R    g0556( .A (n563), .Y (n564) );
  AO21x1_ASAP7_75t_R   g0557( .A1 (n12), .A2 (y2079), .B (x1), .Y (n565) );
  AO21x1_ASAP7_75t_R   g0558( .A1 (n564), .A2 (n565), .B (x4), .Y (n566) );
  AND2x2_ASAP7_75t_R   g0559( .A (n496), .B (n566), .Y (y150) );
  AO21x1_ASAP7_75t_R   g0560( .A1 (y195), .A2 (x4), .B (n539), .Y (y151) );
  AO32x1_ASAP7_75t_R   g0561( .A1 (n352), .A2 (n556), .A3 (x1), .B1 (x0), .B2 (n501), .Y (y152) );
  NAND2x1_ASAP7_75t_R  g0562( .A (n363), .B (n466), .Y (n570) );
  INVx1_ASAP7_75t_R    g0563( .A (n442), .Y (n571) );
  INVx1_ASAP7_75t_R    g0564( .A (n537), .Y (n572) );
  AND3x1_ASAP7_75t_R   g0565( .A (n570), .B (n571), .C (n572), .Y (n573) );
  INVx1_ASAP7_75t_R    g0566( .A (n573), .Y (y153) );
  AO21x1_ASAP7_75t_R   g0567( .A1 (y2079), .A2 (x0), .B (n518), .Y (n575) );
  INVx1_ASAP7_75t_R    g0568( .A (n575), .Y (n576) );
  AO21x1_ASAP7_75t_R   g0569( .A1 (n576), .A2 (x1), .B (n537), .Y (y154) );
  AO21x1_ASAP7_75t_R   g0570( .A1 (n312), .A2 (n497), .B (x4), .Y (n578) );
  AND2x2_ASAP7_75t_R   g0571( .A (n496), .B (n578), .Y (y155) );
  AND2x2_ASAP7_75t_R   g0572( .A (n554), .B (x0), .Y (n580) );
  INVx1_ASAP7_75t_R    g0573( .A (n561), .Y (n581) );
  AO21x1_ASAP7_75t_R   g0574( .A1 (n28), .A2 (n580), .B (n581), .Y (y156) );
  INVx1_ASAP7_75t_R    g0575( .A (n363), .Y (n583) );
  AO21x1_ASAP7_75t_R   g0576( .A1 (y2079), .A2 (x1), .B (x4), .Y (n584) );
  AO21x1_ASAP7_75t_R   g0577( .A1 (n583), .A2 (n16), .B (n584), .Y (n585) );
  INVx1_ASAP7_75t_R    g0578( .A (n585), .Y (n586) );
  AO21x1_ASAP7_75t_R   g0579( .A1 (y195), .A2 (x4), .B (n586), .Y (y157) );
  AO21x1_ASAP7_75t_R   g0580( .A1 (y195), .A2 (x4), .B (n442), .Y (y158) );
  AND3x1_ASAP7_75t_R   g0581( .A (n16), .B (y2079), .C (x0), .Y (n589) );
  AND2x2_ASAP7_75t_R   g0582( .A (n90), .B (y2079), .Y (n590) );
  AO21x1_ASAP7_75t_R   g0583( .A1 (n16), .A2 (x5), .B (x4), .Y (n591) );
  OAI22x1_ASAP7_75t_R  g0584( .A1 (n589), .A2 (n492), .B1 (n590), .B2 (n591), .Y (y159) );
  AO21x1_ASAP7_75t_R   g0585( .A1 (n16), .A2 (n22), .B (y2079), .Y (n593) );
  INVx1_ASAP7_75t_R    g0586( .A (n593), .Y (n594) );
  AO21x1_ASAP7_75t_R   g0587( .A1 (n16), .A2 (x0), .B (n22), .Y (n595) );
  INVx1_ASAP7_75t_R    g0588( .A (n595), .Y (n596) );
  OA21x2_ASAP7_75t_R   g0589( .A1 (n594), .A2 (n596), .B (n387), .Y (y160) );
  AO21x1_ASAP7_75t_R   g0590( .A1 (x5), .A2 (x4), .B (x1), .Y (n598) );
  AO21x1_ASAP7_75t_R   g0591( .A1 (y103), .A2 (n598), .B (n418), .Y (y161) );
  OR3x1_ASAP7_75t_R    g0592( .A (n529), .B (n29), .C (n12), .Y (n600) );
  NAND2x1_ASAP7_75t_R  g0593( .A (n554), .B (n600), .Y (y162) );
  AO21x1_ASAP7_75t_R   g0594( .A1 (n388), .A2 (n28), .B (x1), .Y (n602) );
  AND2x2_ASAP7_75t_R   g0595( .A (n602), .B (y104), .Y (y163) );
  AO21x1_ASAP7_75t_R   g0596( .A1 (y2079), .A2 (x4), .B (x0), .Y (n604) );
  AO21x1_ASAP7_75t_R   g0597( .A1 (x5), .A2 (n22), .B (n604), .Y (n605) );
  INVx1_ASAP7_75t_R    g0598( .A (n598), .Y (n606) );
  AO21x1_ASAP7_75t_R   g0599( .A1 (n12), .A2 (n22), .B (x5), .Y (n607) );
  AND2x2_ASAP7_75t_R   g0600( .A (n28), .B (n607), .Y (n608) );
  OA22x2_ASAP7_75t_R   g0601( .A1 (n605), .A2 (n606), .B1 (n608), .B2 (x1), .Y (y164) );
  AO21x1_ASAP7_75t_R   g0602( .A1 (n15), .A2 (x1), .B (n12), .Y (n610) );
  AO21x1_ASAP7_75t_R   g0603( .A1 (n17), .A2 (x0), .B (n16), .Y (n611) );
  NAND2x1_ASAP7_75t_R  g0604( .A (n610), .B (n611), .Y (y165) );
  AND2x2_ASAP7_75t_R   g0605( .A (n28), .B (n388), .Y (n613) );
  AO21x1_ASAP7_75t_R   g0606( .A1 (n22), .A2 (x0), .B (x5), .Y (n614) );
  NAND2x1_ASAP7_75t_R  g0607( .A (n614), .B (n28), .Y (n615) );
  AO32x1_ASAP7_75t_R   g0608( .A1 (x0), .A2 (n613), .A3 (n312), .B1 (n615), .B2 (x1), .Y (y166) );
  AND2x2_ASAP7_75t_R   g0609( .A (y106), .B (n598), .Y (y167) );
  OR3x1_ASAP7_75t_R    g0610( .A (n337), .B (y2079), .C (x0), .Y (y168) );
  AND3x1_ASAP7_75t_R   g0611( .A (x1), .B (x2), .C (x3), .Y (n619) );
  AO21x1_ASAP7_75t_R   g0612( .A1 (x1), .A2 (x3), .B (x2), .Y (n620) );
  INVx1_ASAP7_75t_R    g0613( .A (n620), .Y (n621) );
  INVx1_ASAP7_75t_R    g0614( .A (n145), .Y (n622) );
  OA33x2_ASAP7_75t_R   g0615( .A1 (x0), .A2 (n619), .A3 (n621), .B1 (n622), .B2 (x2), .B3 (x1), .Y (y169) );
  AO21x1_ASAP7_75t_R   g0616( .A1 (y2079), .A2 (x3), .B (x0), .Y (n624) );
  AO21x1_ASAP7_75t_R   g0617( .A1 (n17), .A2 (n22), .B (n624), .Y (y170) );
  INVx1_ASAP7_75t_R    g0618( .A (n243), .Y (n626) );
  AO21x1_ASAP7_75t_R   g0619( .A1 (n626), .A2 (n241), .B (y69), .Y (y171) );
  INVx1_ASAP7_75t_R    g0620( .A (n316), .Y (n628) );
  OR3x1_ASAP7_75t_R    g0621( .A (x0), .B (x3), .C (x4), .Y (n629) );
  INVx1_ASAP7_75t_R    g0622( .A (n629), .Y (n630) );
  OR3x1_ASAP7_75t_R    g0623( .A (n628), .B (n440), .C (n630), .Y (y172) );
  OR3x1_ASAP7_75t_R    g0624( .A (x3), .B (x4), .C (x5), .Y (n632) );
  AND2x2_ASAP7_75t_R   g0625( .A (y170), .B (n632), .Y (y173) );
  AO21x1_ASAP7_75t_R   g0626( .A1 (n622), .A2 (n128), .B (y69), .Y (y174) );
  AO21x1_ASAP7_75t_R   g0627( .A1 (n377), .A2 (n369), .B (x0), .Y (y175) );
  AO21x1_ASAP7_75t_R   g0628( .A1 (n125), .A2 (y2079), .B (n58), .Y (n636) );
  AO21x1_ASAP7_75t_R   g0629( .A1 (n17), .A2 (n22), .B (n636), .Y (y176) );
  AND3x1_ASAP7_75t_R   g0630( .A (n17), .B (n22), .C (x5), .Y (n638) );
  AO21x1_ASAP7_75t_R   g0631( .A1 (n17), .A2 (n22), .B (x5), .Y (n639) );
  NAND2x1_ASAP7_75t_R  g0632( .A (n12), .B (n639), .Y (n640) );
  AND3x1_ASAP7_75t_R   g0633( .A (n17), .B (y2079), .C (x4), .Y (n641) );
  NAND2x1_ASAP7_75t_R  g0634( .A (x0), .B (n641), .Y (n642) );
  OA21x2_ASAP7_75t_R   g0635( .A1 (n638), .A2 (n640), .B (n642), .Y (y177) );
  AND3x1_ASAP7_75t_R   g0636( .A (n17), .B (y2079), .C (x0), .Y (n644) );
  INVx1_ASAP7_75t_R    g0637( .A (n644), .Y (n645) );
  AND2x2_ASAP7_75t_R   g0638( .A (n645), .B (y168), .Y (y178) );
  AO21x1_ASAP7_75t_R   g0639( .A1 (x4), .A2 (x3), .B (x5), .Y (n647) );
  AO21x1_ASAP7_75t_R   g0640( .A1 (n22), .A2 (n17), .B (n363), .Y (n648) );
  AO21x1_ASAP7_75t_R   g0641( .A1 (x0), .A2 (n647), .B (n648), .Y (y179) );
  AO21x1_ASAP7_75t_R   g0642( .A1 (y2079), .A2 (x3), .B (x4), .Y (n650) );
  INVx1_ASAP7_75t_R    g0643( .A (n650), .Y (n651) );
  AO21x1_ASAP7_75t_R   g0644( .A1 (n22), .A2 (n17), .B (x0), .Y (n652) );
  AND3x1_ASAP7_75t_R   g0645( .A (n382), .B (n652), .C (y2079), .Y (y1828) );
  NOR2x1_ASAP7_75t_R   g0646( .A (n481), .B (y1828), .Y (n654) );
  AO21x1_ASAP7_75t_R   g0647( .A1 (n397), .A2 (n651), .B (n654), .Y (y180) );
  OR3x1_ASAP7_75t_R    g0648( .A (n403), .B (n12), .C (x5), .Y (n656) );
  INVx1_ASAP7_75t_R    g0649( .A (n656), .Y (n657) );
  INVx1_ASAP7_75t_R    g0650( .A (y168), .Y (n658) );
  NOR2x1_ASAP7_75t_R   g0651( .A (n657), .B (n658), .Y (y181) );
  INVx1_ASAP7_75t_R    g0652( .A (n403), .Y (n660) );
  AO21x1_ASAP7_75t_R   g0653( .A1 (n17), .A2 (n22), .B (x0), .Y (n661) );
  AND3x1_ASAP7_75t_R   g0654( .A (n660), .B (n661), .C (y2079), .Y (n662) );
  NOR2x1_ASAP7_75t_R   g0655( .A (n662), .B (n658), .Y (y182) );
  AO21x1_ASAP7_75t_R   g0656( .A1 (n369), .A2 (n290), .B (n58), .Y (y183) );
  AO21x1_ASAP7_75t_R   g0657( .A1 (y2079), .A2 (x2), .B (n544), .Y (n665) );
  AO21x1_ASAP7_75t_R   g0658( .A1 (x0), .A2 (n16), .B (n665), .Y (y184) );
  AO21x1_ASAP7_75t_R   g0659( .A1 (y2079), .A2 (x3), .B (n58), .Y (n667) );
  AO21x1_ASAP7_75t_R   g0660( .A1 (n315), .A2 (n17), .B (n667), .Y (y185) );
  AND3x1_ASAP7_75t_R   g0661( .A (n455), .B (n369), .C (n290), .Y (n669) );
  AO21x1_ASAP7_75t_R   g0662( .A1 (n388), .A2 (x0), .B (n669), .Y (y186) );
  NOR2x1_ASAP7_75t_R   g0663( .A (x3), .B (x5), .Y (n671) );
  INVx1_ASAP7_75t_R    g0664( .A (n671), .Y (n672) );
  OA21x2_ASAP7_75t_R   g0665( .A1 (n529), .A2 (n661), .B (n672), .Y (y187) );
  AO21x1_ASAP7_75t_R   g0666( .A1 (n17), .A2 (n15), .B (n16), .Y (n674) );
  NAND2x1_ASAP7_75t_R  g0667( .A (n12), .B (n674), .Y (y188) );
  NOR2x1_ASAP7_75t_R   g0668( .A (n17), .B (n614), .Y (n676) );
  OR3x1_ASAP7_75t_R    g0669( .A (n676), .B (n58), .C (n337), .Y (y189) );
  AO21x1_ASAP7_75t_R   g0670( .A1 (n17), .A2 (x4), .B (n368), .Y (n678) );
  INVx1_ASAP7_75t_R    g0671( .A (n678), .Y (y2068) );
  AO21x1_ASAP7_75t_R   g0672( .A1 (y2068), .A2 (n310), .B (n58), .Y (y190) );
  OR3x1_ASAP7_75t_R    g0673( .A (x0), .B (x4), .C (x3), .Y (n681) );
  INVx1_ASAP7_75t_R    g0674( .A (n681), .Y (n682) );
  OR3x1_ASAP7_75t_R    g0675( .A (n682), .B (n58), .C (n349), .Y (y191) );
  AO21x1_ASAP7_75t_R   g0676( .A1 (n290), .A2 (n360), .B (x5), .Y (n684) );
  NAND2x1_ASAP7_75t_R  g0677( .A (x5), .B (n328), .Y (n685) );
  INVx1_ASAP7_75t_R    g0678( .A (n330), .Y (n686) );
  AO21x1_ASAP7_75t_R   g0679( .A1 (n684), .A2 (n685), .B (n686), .Y (y192) );
  AO21x1_ASAP7_75t_R   g0680( .A1 (n22), .A2 (n17), .B (y2079), .Y (y3377) );
  AO21x1_ASAP7_75t_R   g0681( .A1 (n382), .A2 (y3377), .B (x0), .Y (y193) );
  AO21x1_ASAP7_75t_R   g0682( .A1 (n16), .A2 (x4), .B (x5), .Y (n690) );
  NAND2x1_ASAP7_75t_R  g0683( .A (n12), .B (n690), .Y (y194) );
  AO21x1_ASAP7_75t_R   g0684( .A1 (n15), .A2 (y2079), .B (n12), .Y (n692) );
  NAND2x1_ASAP7_75t_R  g0685( .A (n692), .B (n312), .Y (y196) );
  AND2x2_ASAP7_75t_R   g0686( .A (n63), .B (n64), .Y (n694) );
  AND2x2_ASAP7_75t_R   g0687( .A (n93), .B (x0), .Y (n695) );
  AO21x1_ASAP7_75t_R   g0688( .A1 (n694), .A2 (n363), .B (n695), .Y (y197) );
  AO21x1_ASAP7_75t_R   g0689( .A1 (n16), .A2 (n22), .B (x5), .Y (n697) );
  AND2x2_ASAP7_75t_R   g0690( .A (n507), .B (y2079), .Y (n698) );
  AO21x1_ASAP7_75t_R   g0691( .A1 (n697), .A2 (x0), .B (n698), .Y (y198) );
  INVx1_ASAP7_75t_R    g0692( .A (n231), .Y (n700) );
  AND3x1_ASAP7_75t_R   g0693( .A (n12), .B (y2079), .C (x2), .Y (n701) );
  AO21x1_ASAP7_75t_R   g0694( .A1 (n700), .A2 (x0), .B (n701), .Y (y200) );
  AO21x1_ASAP7_75t_R   g0695( .A1 (x2), .A2 (x1), .B (n12), .Y (n703) );
  AO21x1_ASAP7_75t_R   g0696( .A1 (n703), .A2 (y2079), .B (n58), .Y (y201) );
  AND3x1_ASAP7_75t_R   g0697( .A (n16), .B (y2079), .C (x2), .Y (n705) );
  INVx1_ASAP7_75t_R    g0698( .A (n705), .Y (n706) );
  AO21x1_ASAP7_75t_R   g0699( .A1 (y2079), .A2 (x2), .B (x0), .Y (n707) );
  AND2x2_ASAP7_75t_R   g0700( .A (n706), .B (n707), .Y (y202) );
  AO21x1_ASAP7_75t_R   g0701( .A1 (n63), .A2 (y2079), .B (x0), .Y (n709) );
  OR3x1_ASAP7_75t_R    g0702( .A (n241), .B (x5), .C (x1), .Y (n710) );
  AND2x2_ASAP7_75t_R   g0703( .A (n709), .B (n710), .Y (y203) );
  AND2x2_ASAP7_75t_R   g0704( .A (n700), .B (n707), .Y (y204) );
  AND3x1_ASAP7_75t_R   g0705( .A (n15), .B (y2079), .C (x0), .Y (n713) );
  INVx1_ASAP7_75t_R    g0706( .A (n713), .Y (n714) );
  AND3x1_ASAP7_75t_R   g0707( .A (n706), .B (n714), .C (y3852), .Y (y205) );
  AND3x1_ASAP7_75t_R   g0708( .A (n63), .B (n64), .C (y2079), .Y (n716) );
  AO21x1_ASAP7_75t_R   g0709( .A1 (x0), .A2 (x5), .B (n716), .Y (y206) );
  AO21x1_ASAP7_75t_R   g0710( .A1 (y2079), .A2 (x0), .B (n22), .Y (n718) );
  NAND2x1_ASAP7_75t_R  g0711( .A (n16), .B (n718), .Y (n719) );
  AND2x2_ASAP7_75t_R   g0712( .A (n719), .B (n387), .Y (y207) );
  AND3x1_ASAP7_75t_R   g0713( .A (n382), .B (n125), .C (y2079), .Y (n721) );
  AO21x1_ASAP7_75t_R   g0714( .A1 (n455), .A2 (x0), .B (n721), .Y (y208) );
  NAND2x1_ASAP7_75t_R  g0715( .A (n12), .B (n647), .Y (y672) );
  OR3x1_ASAP7_75t_R    g0716( .A (x4), .B (x3), .C (x5), .Y (n724) );
  AND2x2_ASAP7_75t_R   g0717( .A (y672), .B (n724), .Y (y209) );
  AO21x1_ASAP7_75t_R   g0718( .A1 (y2079), .A2 (n22), .B (x0), .Y (y1894) );
  OR3x1_ASAP7_75t_R    g0719( .A (x1), .B (x5), .C (x4), .Y (n727) );
  AND2x2_ASAP7_75t_R   g0720( .A (y1894), .B (n727), .Y (y210) );
  OR3x1_ASAP7_75t_R    g0721( .A (y1081), .B (y2079), .C (n109), .Y (y211) );
  AND2x2_ASAP7_75t_R   g0722( .A (n108), .B (y2079), .Y (n730) );
  OR3x1_ASAP7_75t_R    g0723( .A (n730), .B (y1081), .C (n182), .Y (y212) );
  NOR2x1_ASAP7_75t_R   g0724( .A (x2), .B (n488), .Y (n732) );
  OR3x1_ASAP7_75t_R    g0725( .A (n128), .B (y2079), .C (x0), .Y (n733) );
  INVx1_ASAP7_75t_R    g0726( .A (n733), .Y (n734) );
  NOR2x1_ASAP7_75t_R   g0727( .A (n732), .B (n734), .Y (y213) );
  AND3x1_ASAP7_75t_R   g0728( .A (n58), .B (n15), .C (n16), .Y (n736) );
  INVx1_ASAP7_75t_R    g0729( .A (n736), .Y (n737) );
  AO21x1_ASAP7_75t_R   g0730( .A1 (n16), .A2 (n15), .B (y195), .Y (n738) );
  AND2x2_ASAP7_75t_R   g0731( .A (n737), .B (n738), .Y (y214) );
  NAND2x1_ASAP7_75t_R  g0732( .A (x2), .B (y2079), .Y (n740) );
  AO21x1_ASAP7_75t_R   g0733( .A1 (n740), .A2 (n97), .B (n90), .Y (n741) );
  AO21x1_ASAP7_75t_R   g0734( .A1 (n16), .A2 (n15), .B (y2079), .Y (n742) );
  OR3x1_ASAP7_75t_R    g0735( .A (x1), .B (x2), .C (x5), .Y (n743) );
  AO21x1_ASAP7_75t_R   g0736( .A1 (n742), .A2 (n743), .B (x0), .Y (n744) );
  AND2x2_ASAP7_75t_R   g0737( .A (n741), .B (n744), .Y (y215) );
  NAND2x1_ASAP7_75t_R  g0738( .A (x0), .B (n15), .Y (n746) );
  AO21x1_ASAP7_75t_R   g0739( .A1 (n12), .A2 (x2), .B (x1), .Y (n747) );
  AO21x1_ASAP7_75t_R   g0740( .A1 (n746), .A2 (x5), .B (n747), .Y (n748) );
  AND2x2_ASAP7_75t_R   g0741( .A (n748), .B (n733), .Y (y216) );
  AO21x1_ASAP7_75t_R   g0742( .A1 (n16), .A2 (x5), .B (x2), .Y (n750) );
  AO21x1_ASAP7_75t_R   g0743( .A1 (x2), .A2 (x5), .B (x0), .Y (n751) );
  INVx1_ASAP7_75t_R    g0744( .A (n751), .Y (n752) );
  AO21x1_ASAP7_75t_R   g0745( .A1 (x2), .A2 (x5), .B (x1), .Y (n753) );
  AND2x2_ASAP7_75t_R   g0746( .A (n753), .B (x0), .Y (n754) );
  AO21x1_ASAP7_75t_R   g0747( .A1 (n750), .A2 (n752), .B (n754), .Y (y217) );
  AND2x2_ASAP7_75t_R   g0748( .A (x2), .B (x5), .Y (n756) );
  INVx1_ASAP7_75t_R    g0749( .A (n756), .Y (n757) );
  AO21x1_ASAP7_75t_R   g0750( .A1 (n15), .A2 (y2079), .B (n16), .Y (n758) );
  AND3x1_ASAP7_75t_R   g0751( .A (n757), .B (n758), .C (x0), .Y (n759) );
  NOR2x1_ASAP7_75t_R   g0752( .A (n759), .B (n734), .Y (y218) );
  AND3x1_ASAP7_75t_R   g0753( .A (n15), .B (n16), .C (x0), .Y (n761) );
  INVx1_ASAP7_75t_R    g0754( .A (n761), .Y (n762) );
  AO21x1_ASAP7_75t_R   g0755( .A1 (x2), .A2 (x1), .B (x5), .Y (n763) );
  AO32x1_ASAP7_75t_R   g0756( .A1 (n67), .A2 (n762), .A3 (n763), .B1 (n52), .B2 (n363), .Y (y219) );
  INVx1_ASAP7_75t_R    g0757( .A (n58), .Y (n765) );
  AND2x2_ASAP7_75t_R   g0758( .A (y3852), .B (n753), .Y (y3732) );
  AO21x1_ASAP7_75t_R   g0759( .A1 (n765), .A2 (n128), .B (y3732), .Y (y220) );
  AND2x2_ASAP7_75t_R   g0760( .A (n707), .B (n753), .Y (y555) );
  AO21x1_ASAP7_75t_R   g0761( .A1 (n765), .A2 (n128), .B (y555), .Y (y221) );
  AO21x1_ASAP7_75t_R   g0762( .A1 (n740), .A2 (n97), .B (x1), .Y (n770) );
  INVx1_ASAP7_75t_R    g0763( .A (n770), .Y (n771) );
  AND3x1_ASAP7_75t_R   g0764( .A (n15), .B (x5), .C (x0), .Y (n772) );
  AO21x1_ASAP7_75t_R   g0765( .A1 (y2079), .A2 (x2), .B (n772), .Y (n773) );
  INVx1_ASAP7_75t_R    g0766( .A (n773), .Y (n774) );
  OA22x2_ASAP7_75t_R   g0767( .A1 (n707), .A2 (n771), .B1 (n774), .B2 (x1), .Y (y222) );
  INVx1_ASAP7_75t_R    g0768( .A (n544), .Y (n776) );
  AO21x1_ASAP7_75t_R   g0769( .A1 (n776), .A2 (n64), .B (n58), .Y (n777) );
  AO21x1_ASAP7_75t_R   g0770( .A1 (n312), .A2 (n497), .B (n746), .Y (n778) );
  AND2x2_ASAP7_75t_R   g0771( .A (n777), .B (n778), .Y (y223) );
  INVx1_ASAP7_75t_R    g0772( .A (n753), .Y (n780) );
  AO21x1_ASAP7_75t_R   g0773( .A1 (y2079), .A2 (x0), .B (n16), .Y (n781) );
  NAND2x1_ASAP7_75t_R  g0774( .A (n15), .B (n781), .Y (n782) );
  AO32x1_ASAP7_75t_R   g0775( .A1 (n583), .A2 (n692), .A3 (n780), .B1 (y2389), .B2 (n782), .Y (y224) );
  OR3x1_ASAP7_75t_R    g0776( .A (n544), .B (n12), .C (x2), .Y (n784) );
  AND2x2_ASAP7_75t_R   g0777( .A (n777), .B (n784), .Y (y225) );
  AND3x1_ASAP7_75t_R   g0778( .A (n733), .B (n784), .C (n700), .Y (y226) );
  AND3x1_ASAP7_75t_R   g0779( .A (y2079), .B (x1), .C (x2), .Y (n787) );
  OR3x1_ASAP7_75t_R    g0780( .A (n787), .B (n58), .C (n51), .Y (n788) );
  AND2x2_ASAP7_75t_R   g0781( .A (n788), .B (n762), .Y (y227) );
  AND2x2_ASAP7_75t_R   g0782( .A (n757), .B (n758), .Y (n790) );
  AND3x1_ASAP7_75t_R   g0783( .A (n128), .B (n12), .C (x5), .Y (n791) );
  INVx1_ASAP7_75t_R    g0784( .A (n791), .Y (n792) );
  OAI21x1_ASAP7_75t_R  g0785( .A1 (n481), .A2 (n790), .B (n792), .Y (y228) );
  AO21x1_ASAP7_75t_R   g0786( .A1 (n312), .A2 (n497), .B (x2), .Y (n794) );
  INVx1_ASAP7_75t_R    g0787( .A (n794), .Y (n795) );
  OA21x2_ASAP7_75t_R   g0788( .A1 (n795), .A2 (x0), .B (n737), .Y (y229) );
  AO21x1_ASAP7_75t_R   g0789( .A1 (n16), .A2 (n15), .B (n12), .Y (n797) );
  INVx1_ASAP7_75t_R    g0790( .A (n797), .Y (n798) );
  AO21x1_ASAP7_75t_R   g0791( .A1 (n776), .A2 (n241), .B (n798), .Y (y230) );
  AO21x1_ASAP7_75t_R   g0792( .A1 (x1), .A2 (x5), .B (x2), .Y (n800) );
  INVx1_ASAP7_75t_R    g0793( .A (n800), .Y (n801) );
  INVx1_ASAP7_75t_R    g0794( .A (n732), .Y (n802) );
  OA21x2_ASAP7_75t_R   g0795( .A1 (x0), .A2 (n801), .B (n802), .Y (y231) );
  NAND2x1_ASAP7_75t_R  g0796( .A (n108), .B (n155), .Y (y232) );
  AO21x1_ASAP7_75t_R   g0797( .A1 (n77), .A2 (n674), .B (x0), .Y (n805) );
  OR3x1_ASAP7_75t_R    g0798( .A (n76), .B (n12), .C (x1), .Y (n806) );
  AND2x2_ASAP7_75t_R   g0799( .A (n805), .B (n806), .Y (y233) );
  AO21x1_ASAP7_75t_R   g0800( .A1 (n137), .A2 (n72), .B (n90), .Y (n808) );
  AO21x1_ASAP7_75t_R   g0801( .A1 (x2), .A2 (x3), .B (x1), .Y (n809) );
  NAND2x1_ASAP7_75t_R  g0802( .A (n12), .B (n809), .Y (n810) );
  AND2x2_ASAP7_75t_R   g0803( .A (n808), .B (n810), .Y (y234) );
  INVx1_ASAP7_75t_R    g0804( .A (n213), .Y (n812) );
  AND2x2_ASAP7_75t_R   g0805( .A (n809), .B (x0), .Y (n813) );
  AO21x1_ASAP7_75t_R   g0806( .A1 (n812), .A2 (n16), .B (n813), .Y (y235) );
  AND2x2_ASAP7_75t_R   g0807( .A (n397), .B (x4), .Y (n815) );
  AO21x1_ASAP7_75t_R   g0808( .A1 (n341), .A2 (x3), .B (n815), .Y (y236) );
  AND3x1_ASAP7_75t_R   g0809( .A (n14), .B (n18), .C (x0), .Y (n817) );
  INVx1_ASAP7_75t_R    g0810( .A (n817), .Y (n818) );
  AO21x1_ASAP7_75t_R   g0811( .A1 (n14), .A2 (n18), .B (x0), .Y (n819) );
  AND2x2_ASAP7_75t_R   g0812( .A (n818), .B (n819), .Y (y237) );
  NAND2x1_ASAP7_75t_R  g0813( .A (x5), .B (n155), .Y (y238) );
  AO21x1_ASAP7_75t_R   g0814( .A1 (n129), .A2 (x0), .B (n363), .Y (y239) );
  AND2x2_ASAP7_75t_R   g0815( .A (n129), .B (y3852), .Y (y240) );
  AO21x1_ASAP7_75t_R   g0816( .A1 (n16), .A2 (x2), .B (x5), .Y (n824) );
  NAND2x1_ASAP7_75t_R  g0817( .A (n12), .B (n824), .Y (n825) );
  AND3x1_ASAP7_75t_R   g0818( .A (n16), .B (n15), .C (x0), .Y (n826) );
  INVx1_ASAP7_75t_R    g0819( .A (n826), .Y (n827) );
  AND2x2_ASAP7_75t_R   g0820( .A (n825), .B (n827), .Y (y241) );
  NAND2x1_ASAP7_75t_R  g0821( .A (n797), .B (n312), .Y (y242) );
  INVx1_ASAP7_75t_R    g0822( .A (n716), .Y (n830) );
  NAND2x1_ASAP7_75t_R  g0823( .A (n12), .B (n830), .Y (y1714) );
  AND2x2_ASAP7_75t_R   g0824( .A (y1714), .B (n762), .Y (y243) );
  OR3x1_ASAP7_75t_R    g0825( .A (n756), .B (n12), .C (x1), .Y (n833) );
  AND2x2_ASAP7_75t_R   g0826( .A (n833), .B (y3852), .Y (y244) );
  AO21x1_ASAP7_75t_R   g0827( .A1 (y2079), .A2 (x0), .B (n15), .Y (n835) );
  NAND2x1_ASAP7_75t_R  g0828( .A (n16), .B (n835), .Y (n836) );
  AND2x2_ASAP7_75t_R   g0829( .A (n836), .B (y3852), .Y (y245) );
  AO21x1_ASAP7_75t_R   g0830( .A1 (n700), .A2 (x0), .B (n363), .Y (n838) );
  AND3x1_ASAP7_75t_R   g0831( .A (n231), .B (n15), .C (x0), .Y (n839) );
  AO21x1_ASAP7_75t_R   g0832( .A1 (n838), .A2 (n782), .B (n839), .Y (y246) );
  AO21x1_ASAP7_75t_R   g0833( .A1 (n16), .A2 (y2079), .B (n15), .Y (n841) );
  AO21x1_ASAP7_75t_R   g0834( .A1 (n776), .A2 (n841), .B (n12), .Y (n842) );
  NAND2x1_ASAP7_75t_R  g0835( .A (n583), .B (n842), .Y (y247) );
  AO21x1_ASAP7_75t_R   g0836( .A1 (n740), .A2 (n746), .B (x1), .Y (n844) );
  AND2x2_ASAP7_75t_R   g0837( .A (n844), .B (n709), .Y (y248) );
  AO21x1_ASAP7_75t_R   g0838( .A1 (n746), .A2 (x1), .B (n826), .Y (n846) );
  OR3x1_ASAP7_75t_R    g0839( .A (n128), .B (y2079), .C (n12), .Y (n847) );
  INVx1_ASAP7_75t_R    g0840( .A (n847), .Y (n848) );
  AO21x1_ASAP7_75t_R   g0841( .A1 (y2079), .A2 (n846), .B (n848), .Y (y249) );
  AND2x2_ASAP7_75t_R   g0842( .A (n782), .B (y2389), .Y (y251) );
  AO21x1_ASAP7_75t_R   g0843( .A1 (n15), .A2 (x0), .B (x1), .Y (n851) );
  AO32x1_ASAP7_75t_R   g0844( .A1 (y2079), .A2 (n63), .A3 (n851), .B1 (n58), .B2 (n129), .Y (y252) );
  NAND2x1_ASAP7_75t_R  g0845( .A (n763), .B (n155), .Y (y253) );
  NOR2x1_ASAP7_75t_R   g0846( .A (x5), .B (y25), .Y (n854) );
  AO21x1_ASAP7_75t_R   g0847( .A1 (n52), .A2 (x0), .B (n854), .Y (y254) );
  NOR2x1_ASAP7_75t_R   g0848( .A (x2), .B (x5), .Y (n856) );
  AO21x1_ASAP7_75t_R   g0849( .A1 (n129), .A2 (x0), .B (n856), .Y (y255) );
  AO21x1_ASAP7_75t_R   g0850( .A1 (n15), .A2 (y2079), .B (x0), .Y (n858) );
  AND2x2_ASAP7_75t_R   g0851( .A (n827), .B (n858), .Y (y256) );
  NAND2x1_ASAP7_75t_R  g0852( .A (n17), .B (n56), .Y (n860) );
  INVx1_ASAP7_75t_R    g0853( .A (n860), .Y (n861) );
  OA21x2_ASAP7_75t_R   g0854( .A1 (n861), .A2 (n141), .B (n238), .Y (y257) );
  AO21x1_ASAP7_75t_R   g0855( .A1 (n17), .A2 (x0), .B (n15), .Y (n863) );
  NAND2x1_ASAP7_75t_R  g0856( .A (n16), .B (n863), .Y (n864) );
  AO21x1_ASAP7_75t_R   g0857( .A1 (x1), .A2 (x2), .B (x3), .Y (n865) );
  NAND2x1_ASAP7_75t_R  g0858( .A (n12), .B (n865), .Y (n866) );
  AND2x2_ASAP7_75t_R   g0859( .A (n864), .B (n866), .Y (y258) );
  AO21x1_ASAP7_75t_R   g0860( .A1 (n137), .A2 (n72), .B (x1), .Y (n868) );
  NAND2x1_ASAP7_75t_R  g0861( .A (n12), .B (n117), .Y (n869) );
  INVx1_ASAP7_75t_R    g0862( .A (n869), .Y (n870) );
  AO21x1_ASAP7_75t_R   g0863( .A1 (n868), .A2 (x0), .B (n870), .Y (y259) );
  OR3x1_ASAP7_75t_R    g0864( .A (n211), .B (n12), .C (x1), .Y (n872) );
  AND2x2_ASAP7_75t_R   g0865( .A (n872), .B (n116), .Y (y260) );
  AO21x1_ASAP7_75t_R   g0866( .A1 (n16), .A2 (n17), .B (n15), .Y (n874) );
  AO21x1_ASAP7_75t_R   g0867( .A1 (n626), .A2 (n874), .B (n12), .Y (n875) );
  INVx1_ASAP7_75t_R    g0868( .A (n158), .Y (n876) );
  NAND2x1_ASAP7_75t_R  g0869( .A (n875), .B (n876), .Y (y261) );
  AO21x1_ASAP7_75t_R   g0870( .A1 (x2), .A2 (x1), .B (x3), .Y (n878) );
  NAND2x1_ASAP7_75t_R  g0871( .A (x0), .B (n878), .Y (n879) );
  INVx1_ASAP7_75t_R    g0872( .A (n879), .Y (n880) );
  OA21x2_ASAP7_75t_R   g0873( .A1 (n158), .A2 (n880), .B (n52), .Y (y262) );
  AO21x1_ASAP7_75t_R   g0874( .A1 (n809), .A2 (x0), .B (n45), .Y (y263) );
  AO21x1_ASAP7_75t_R   g0875( .A1 (x3), .A2 (x2), .B (x1), .Y (n883) );
  AND2x2_ASAP7_75t_R   g0876( .A (n883), .B (x0), .Y (y2826) );
  AO21x1_ASAP7_75t_R   g0877( .A1 (y9), .A2 (n81), .B (y2826), .Y (y264) );
  AO21x1_ASAP7_75t_R   g0878( .A1 (n137), .A2 (n746), .B (x1), .Y (n886) );
  AND2x2_ASAP7_75t_R   g0879( .A (n886), .B (n116), .Y (y265) );
  AO21x1_ASAP7_75t_R   g0880( .A1 (n661), .A2 (x5), .B (n676), .Y (y266) );
  NOR2x1_ASAP7_75t_R   g0881( .A (n12), .B (n128), .Y (n889) );
  INVx1_ASAP7_75t_R    g0882( .A (n865), .Y (n890) );
  AO21x1_ASAP7_75t_R   g0883( .A1 (n63), .A2 (n64), .B (n125), .Y (n891) );
  OA211x2_ASAP7_75t_R  g0884( .A1 (n889), .A2 (n890), .B (n891), .C (y9), .Y (y267) );
  AND2x2_ASAP7_75t_R   g0885( .A (n169), .B (n883), .Y (y268) );
  NOR2x1_ASAP7_75t_R   g0886( .A (n12), .B (n20), .Y (y269) );
  OR3x1_ASAP7_75t_R    g0887( .A (x3), .B (x2), .C (x1), .Y (n895) );
  INVx1_ASAP7_75t_R    g0888( .A (n895), .Y (n896) );
  OR3x1_ASAP7_75t_R    g0889( .A (n13), .B (n12), .C (x3), .Y (n897) );
  OA21x2_ASAP7_75t_R   g0890( .A1 (y1081), .A2 (n896), .B (n897), .Y (y270) );
  AO21x1_ASAP7_75t_R   g0891( .A1 (n90), .A2 (n219), .B (n22), .Y (n899) );
  NOR2x1_ASAP7_75t_R   g0892( .A (y2079), .B (n899), .Y (n900) );
  INVx1_ASAP7_75t_R    g0893( .A (n900), .Y (y271) );
  AO21x1_ASAP7_75t_R   g0894( .A1 (n219), .A2 (n90), .B (n22), .Y (n902) );
  NOR2x1_ASAP7_75t_R   g0895( .A (y2079), .B (n902), .Y (n903) );
  NOR2x1_ASAP7_75t_R   g0896( .A (n532), .B (n903), .Y (y272) );
  AND3x1_ASAP7_75t_R   g0897( .A (n90), .B (n219), .C (n22), .Y (n905) );
  NAND2x1_ASAP7_75t_R  g0898( .A (y2079), .B (n905), .Y (n906) );
  AND2x2_ASAP7_75t_R   g0899( .A (y271), .B (n906), .Y (y273) );
  AO21x1_ASAP7_75t_R   g0900( .A1 (n219), .A2 (n90), .B (y2079), .Y (n908) );
  AO21x1_ASAP7_75t_R   g0901( .A1 (n908), .A2 (n490), .B (n29), .Y (y274) );
  AO21x1_ASAP7_75t_R   g0902( .A1 (x1), .A2 (x0), .B (n22), .Y (n910) );
  AND2x2_ASAP7_75t_R   g0903( .A (n910), .B (x5), .Y (n911) );
  OR3x1_ASAP7_75t_R    g0904( .A (n911), .B (n227), .C (n529), .Y (y275) );
  AO21x1_ASAP7_75t_R   g0905( .A1 (n12), .A2 (n16), .B (y2079), .Y (n913) );
  INVx1_ASAP7_75t_R    g0906( .A (n310), .Y (n914) );
  AO221x2_ASAP7_75t_R  g0907( .A1 (n913), .A2 (n501), .B1 (n299), .B2 (n544), .C (n914), .Y (y276) );
  AO21x1_ASAP7_75t_R   g0908( .A1 (x1), .A2 (x5), .B (n22), .Y (n916) );
  NAND2x1_ASAP7_75t_R  g0909( .A (n12), .B (n916), .Y (n917) );
  AND3x1_ASAP7_75t_R   g0910( .A (n537), .B (n16), .C (x5), .Y (n918) );
  INVx1_ASAP7_75t_R    g0911( .A (n918), .Y (n919) );
  OA21x2_ASAP7_75t_R   g0912( .A1 (n442), .A2 (n917), .B (n919), .Y (y277) );
  AND3x1_ASAP7_75t_R   g0913( .A (n556), .B (n352), .C (n17), .Y (n921) );
  NAND2x1_ASAP7_75t_R  g0914( .A (x3), .B (n386), .Y (n922) );
  INVx1_ASAP7_75t_R    g0915( .A (n922), .Y (n923) );
  NOR2x1_ASAP7_75t_R   g0916( .A (n921), .B (n923), .Y (y278) );
  INVx1_ASAP7_75t_R    g0917( .A (n9), .Y (n925) );
  AO21x1_ASAP7_75t_R   g0918( .A1 (n14), .A2 (n18), .B (n12), .Y (n926) );
  NAND2x1_ASAP7_75t_R  g0919( .A (n895), .B (n926), .Y (y514) );
  AO21x1_ASAP7_75t_R   g0920( .A1 (n925), .A2 (n674), .B (y514), .Y (y279) );
  NOR2x1_ASAP7_75t_R   g0921( .A (x1), .B (n429), .Y (n929) );
  INVx1_ASAP7_75t_R    g0922( .A (n929), .Y (n930) );
  OR3x1_ASAP7_75t_R    g0923( .A (n43), .B (n22), .C (y2079), .Y (n931) );
  AO21x1_ASAP7_75t_R   g0924( .A1 (n930), .A2 (n931), .B (n143), .Y (y280) );
  NOR2x1_ASAP7_75t_R   g0925( .A (n839), .B (n481), .Y (y281) );
  AO21x1_ASAP7_75t_R   g0926( .A1 (x5), .A2 (x4), .B (n12), .Y (n934) );
  AO21x1_ASAP7_75t_R   g0927( .A1 (y103), .A2 (n419), .B (n16), .Y (n935) );
  OAI21x1_ASAP7_75t_R  g0928( .A1 (n410), .A2 (n457), .B (n935), .Y (n936) );
  NAND2x1_ASAP7_75t_R  g0929( .A (n934), .B (n936), .Y (y282) );
  AO21x1_ASAP7_75t_R   g0930( .A1 (x1), .A2 (x4), .B (x0), .Y (n938) );
  AND2x2_ASAP7_75t_R   g0931( .A (n436), .B (n466), .Y (n939) );
  INVx1_ASAP7_75t_R    g0932( .A (n939), .Y (n940) );
  AO221x2_ASAP7_75t_R  g0933( .A1 (n593), .A2 (n938), .B1 (n481), .B2 (n940), .C (n143), .Y (y283) );
  AO21x1_ASAP7_75t_R   g0934( .A1 (n90), .A2 (n219), .B (y2079), .Y (y1873) );
  NOR2x1_ASAP7_75t_R   g0935( .A (n22), .B (y1873), .Y (n943) );
  AND3x1_ASAP7_75t_R   g0936( .A (y3293), .B (n90), .C (n219), .Y (y1635) );
  AND2x2_ASAP7_75t_R   g0937( .A (y1635), .B (n523), .Y (n945) );
  NOR2x1_ASAP7_75t_R   g0938( .A (n943), .B (n945), .Y (y284) );
  OR3x1_ASAP7_75t_R    g0939( .A (x1), .B (x0), .C (x4), .Y (n947) );
  AO21x1_ASAP7_75t_R   g0940( .A1 (n16), .A2 (n12), .B (n22), .Y (n948) );
  NAND2x1_ASAP7_75t_R  g0941( .A (n947), .B (n948), .Y (n949) );
  AND3x1_ASAP7_75t_R   g0942( .A (n16), .B (n12), .C (x4), .Y (n950) );
  AO21x1_ASAP7_75t_R   g0943( .A1 (n466), .A2 (x0), .B (n950), .Y (n951) );
  OA22x2_ASAP7_75t_R   g0944( .A1 (n949), .A2 (x5), .B1 (n951), .B2 (n463), .Y (y285) );
  AO21x1_ASAP7_75t_R   g0945( .A1 (n228), .A2 (y3293), .B (y863), .Y (n953) );
  NAND2x1_ASAP7_75t_R  g0946( .A (x5), .B (n950), .Y (y3234) );
  INVx1_ASAP7_75t_R    g0947( .A (y3234), .Y (n955) );
  AO21x1_ASAP7_75t_R   g0948( .A1 (n419), .A2 (n953), .B (n955), .Y (y286) );
  AO21x1_ASAP7_75t_R   g0949( .A1 (y2079), .A2 (x4), .B (n143), .Y (n957) );
  AO21x1_ASAP7_75t_R   g0950( .A1 (n16), .A2 (n307), .B (n957), .Y (y287) );
  AND3x1_ASAP7_75t_R   g0951( .A (y2079), .B (n22), .C (x3), .Y (n959) );
  NOR2x1_ASAP7_75t_R   g0952( .A (n410), .B (n959), .Y (y288) );
  AO21x1_ASAP7_75t_R   g0953( .A1 (n16), .A2 (x4), .B (y2079), .Y (n961) );
  INVx1_ASAP7_75t_R    g0954( .A (n961), .Y (n962) );
  AO21x1_ASAP7_75t_R   g0955( .A1 (y2079), .A2 (n436), .B (n962), .Y (n963) );
  AO21x1_ASAP7_75t_R   g0956( .A1 (x1), .A2 (x5), .B (x0), .Y (n964) );
  INVx1_ASAP7_75t_R    g0957( .A (n964), .Y (n965) );
  AO21x1_ASAP7_75t_R   g0958( .A1 (n963), .A2 (x0), .B (n965), .Y (y289) );
  AND3x1_ASAP7_75t_R   g0959( .A (n16), .B (x4), .C (x0), .Y (n967) );
  INVx1_ASAP7_75t_R    g0960( .A (n967), .Y (n968) );
  AO21x1_ASAP7_75t_R   g0961( .A1 (n12), .A2 (x1), .B (y2079), .Y (n969) );
  INVx1_ASAP7_75t_R    g0962( .A (n969), .Y (n970) );
  AO21x1_ASAP7_75t_R   g0963( .A1 (n12), .A2 (x1), .B (x4), .Y (n971) );
  AND2x2_ASAP7_75t_R   g0964( .A (n971), .B (y2079), .Y (n972) );
  AO21x1_ASAP7_75t_R   g0965( .A1 (n968), .A2 (n970), .B (n972), .Y (y290) );
  AND3x1_ASAP7_75t_R   g0966( .A (n12), .B (n16), .C (x4), .Y (n974) );
  NOR2x1_ASAP7_75t_R   g0967( .A (x5), .B (n974), .Y (n975) );
  AO21x1_ASAP7_75t_R   g0968( .A1 (n16), .A2 (x4), .B (n12), .Y (n976) );
  INVx1_ASAP7_75t_R    g0969( .A (n976), .Y (n977) );
  AND3x1_ASAP7_75t_R   g0970( .A (n12), .B (n16), .C (x5), .Y (n978) );
  OR3x1_ASAP7_75t_R    g0971( .A (n975), .B (n977), .C (n978), .Y (y291) );
  NAND2x1_ASAP7_75t_R  g0972( .A (n527), .B (n352), .Y (n980) );
  INVx1_ASAP7_75t_R    g0973( .A (n980), .Y (n981) );
  AO21x1_ASAP7_75t_R   g0974( .A1 (y3852), .A2 (x1), .B (n978), .Y (n982) );
  OR3x1_ASAP7_75t_R    g0975( .A (n527), .B (n12), .C (x5), .Y (n983) );
  INVx1_ASAP7_75t_R    g0976( .A (n983), .Y (n984) );
  OR3x1_ASAP7_75t_R    g0977( .A (n981), .B (n982), .C (n984), .Y (y292) );
  AND2x2_ASAP7_75t_R   g0978( .A (n129), .B (n858), .Y (y293) );
  NOR2x1_ASAP7_75t_R   g0979( .A (n537), .B (n497), .Y (n987) );
  AO21x1_ASAP7_75t_R   g0980( .A1 (n12), .A2 (x5), .B (n16), .Y (n988) );
  INVx1_ASAP7_75t_R    g0981( .A (n988), .Y (n989) );
  AND3x1_ASAP7_75t_R   g0982( .A (y2079), .B (x4), .C (x0), .Y (n990) );
  OR3x1_ASAP7_75t_R    g0983( .A (n987), .B (n989), .C (n990), .Y (y294) );
  NOR2x1_ASAP7_75t_R   g0984( .A (n12), .B (n53), .Y (y295) );
  INVx1_ASAP7_75t_R    g0985( .A (n497), .Y (n993) );
  AO21x1_ASAP7_75t_R   g0986( .A1 (y2079), .A2 (x0), .B (x1), .Y (n994) );
  AND2x2_ASAP7_75t_R   g0987( .A (n604), .B (n994), .Y (n995) );
  AO21x1_ASAP7_75t_R   g0988( .A1 (n572), .A2 (n993), .B (n995), .Y (y296) );
  AND2x2_ASAP7_75t_R   g0989( .A (n312), .B (n497), .Y (n997) );
  INVx1_ASAP7_75t_R    g0990( .A (n997), .Y (n998) );
  AND2x2_ASAP7_75t_R   g0991( .A (x1), .B (x4), .Y (n999) );
  AO21x1_ASAP7_75t_R   g0992( .A1 (n22), .A2 (x5), .B (n999), .Y (n1000) );
  OR3x1_ASAP7_75t_R    g0993( .A (n1000), .B (n12), .C (n231), .Y (n1001) );
  OA21x2_ASAP7_75t_R   g0994( .A1 (n998), .A2 (x0), .B (n1001), .Y (y297) );
  AND3x1_ASAP7_75t_R   g0995( .A (n219), .B (n90), .C (x5), .Y (n1003) );
  NOR2x1_ASAP7_75t_R   g0996( .A (n43), .B (n388), .Y (n1004) );
  OR3x1_ASAP7_75t_R    g0997( .A (n1003), .B (n1004), .C (n527), .Y (y298) );
  AO21x1_ASAP7_75t_R   g0998( .A1 (n968), .A2 (n219), .B (y2079), .Y (y2442) );
  AO21x1_ASAP7_75t_R   g0999( .A1 (n12), .A2 (n16), .B (n22), .Y (n1007) );
  NAND2x1_ASAP7_75t_R  g1000( .A (y2079), .B (n1007), .Y (n1008) );
  AND2x2_ASAP7_75t_R   g1001( .A (y2442), .B (n1008), .Y (y299) );
  OR3x1_ASAP7_75t_R    g1002( .A (n982), .B (n977), .C (n974), .Y (y300) );
  AO21x1_ASAP7_75t_R   g1003( .A1 (y2079), .A2 (x4), .B (n16), .Y (n1011) );
  NOR2x1_ASAP7_75t_R   g1004( .A (x0), .B (n1011), .Y (n1012) );
  NOR2x1_ASAP7_75t_R   g1005( .A (n967), .B (n1012), .Y (y301) );
  AO21x1_ASAP7_75t_R   g1006( .A1 (n455), .A2 (n965), .B (n977), .Y (y302) );
  AO32x1_ASAP7_75t_R   g1007( .A1 (n776), .A2 (n455), .A3 (n572), .B1 (x1), .B2 (x0), .Y (y303) );
  AND3x1_ASAP7_75t_R   g1008( .A (y3852), .B (n352), .C (x1), .Y (n1016) );
  AND3x1_ASAP7_75t_R   g1009( .A (x0), .B (x1), .C (x4), .Y (n1017) );
  OR3x1_ASAP7_75t_R    g1010( .A (n1016), .B (n1017), .C (n512), .Y (y304) );
  AO21x1_ASAP7_75t_R   g1011( .A1 (n22), .A2 (n17), .B (n374), .Y (n1019) );
  INVx1_ASAP7_75t_R    g1012( .A (n1019), .Y (n1020) );
  OA21x2_ASAP7_75t_R   g1013( .A1 (n1020), .A2 (n363), .B (n684), .Y (y305) );
  AND3x1_ASAP7_75t_R   g1014( .A (n219), .B (n90), .C (n22), .Y (n1022) );
  NAND2x1_ASAP7_75t_R  g1015( .A (y2079), .B (n1022), .Y (n1023) );
  NAND2x1_ASAP7_75t_R  g1016( .A (n511), .B (n988), .Y (y630) );
  AND2x2_ASAP7_75t_R   g1017( .A (n1023), .B (y630), .Y (y306) );
  OR3x1_ASAP7_75t_R    g1018( .A (n16), .B (y2079), .C (x0), .Y (n1026) );
  NAND2x1_ASAP7_75t_R  g1019( .A (n90), .B (n1026), .Y (n1027) );
  INVx1_ASAP7_75t_R    g1020( .A (n1027), .Y (n1028) );
  AND3x1_ASAP7_75t_R   g1021( .A (n16), .B (n22), .C (x0), .Y (n1029) );
  AO21x1_ASAP7_75t_R   g1022( .A1 (n1028), .A2 (n455), .B (n1029), .Y (y307) );
  AO21x1_ASAP7_75t_R   g1023( .A1 (n1000), .A2 (y3852), .B (n43), .Y (y308) );
  INVx1_ASAP7_75t_R    g1024( .A (n84), .Y (n1032) );
  AND3x1_ASAP7_75t_R   g1025( .A (n15), .B (n16), .C (x3), .Y (n1033) );
  NOR2x1_ASAP7_75t_R   g1026( .A (n12), .B (n1033), .Y (n1034) );
  AO21x1_ASAP7_75t_R   g1027( .A1 (n694), .A2 (n1032), .B (n1034), .Y (y309) );
  AO21x1_ASAP7_75t_R   g1028( .A1 (n12), .A2 (x4), .B (x5), .Y (n1036) );
  INVx1_ASAP7_75t_R    g1029( .A (n1036), .Y (y2147) );
  AO21x1_ASAP7_75t_R   g1030( .A1 (n968), .A2 (n219), .B (y2147), .Y (y310) );
  NAND2x1_ASAP7_75t_R  g1031( .A (n16), .B (y1894), .Y (n1039) );
  OR3x1_ASAP7_75t_R    g1032( .A (n418), .B (n16), .C (x0), .Y (n1040) );
  INVx1_ASAP7_75t_R    g1033( .A (n934), .Y (y1378) );
  AO21x1_ASAP7_75t_R   g1034( .A1 (n1039), .A2 (n1040), .B (y1378), .Y (y311) );
  AND3x1_ASAP7_75t_R   g1035( .A (n672), .B (n556), .C (n360), .Y (y2723) );
  OR2x4_ASAP7_75t_R    g1036( .A (x0), .B (y2723), .Y (y312) );
  AND3x1_ASAP7_75t_R   g1037( .A (n388), .B (n28), .C (n16), .Y (n1045) );
  INVx1_ASAP7_75t_R    g1038( .A (n1045), .Y (n1046) );
  AO21x1_ASAP7_75t_R   g1039( .A1 (n22), .A2 (y2079), .B (x0), .Y (n1047) );
  AO21x1_ASAP7_75t_R   g1040( .A1 (n1046), .A2 (n1047), .B (n43), .Y (y313) );
  OR3x1_ASAP7_75t_R    g1041( .A (y772), .B (n478), .C (n974), .Y (y314) );
  AO21x1_ASAP7_75t_R   g1042( .A1 (n22), .A2 (y2079), .B (n16), .Y (n1050) );
  INVx1_ASAP7_75t_R    g1043( .A (n513), .Y (n1051) );
  AO21x1_ASAP7_75t_R   g1044( .A1 (n455), .A2 (n143), .B (n1051), .Y (y621) );
  AO21x1_ASAP7_75t_R   g1045( .A1 (n12), .A2 (n1050), .B (y621), .Y (y315) );
  AND3x1_ASAP7_75t_R   g1046( .A (n90), .B (y2079), .C (n22), .Y (n1054) );
  NAND2x1_ASAP7_75t_R  g1047( .A (n511), .B (n180), .Y (y3274) );
  XOR2x2_ASAP7_75t_R   g1048( .A (n1054), .B (y3274), .Y (y316) );
  OA21x2_ASAP7_75t_R   g1049( .A1 (n29), .A2 (n31), .B (x0), .Y (y689) );
  AO21x1_ASAP7_75t_R   g1050( .A1 (n12), .A2 (n523), .B (y689), .Y (y317) );
  AO21x1_ASAP7_75t_R   g1051( .A1 (x0), .A2 (x5), .B (x1), .Y (n1059) );
  INVx1_ASAP7_75t_R    g1052( .A (n1059), .Y (n1060) );
  AO21x1_ASAP7_75t_R   g1053( .A1 (n1000), .A2 (x0), .B (n1060), .Y (y318) );
  INVx1_ASAP7_75t_R    g1054( .A (n45), .Y (n1062) );
  AO21x1_ASAP7_75t_R   g1055( .A1 (n228), .A2 (n1062), .B (n216), .Y (y319) );
  INVx1_ASAP7_75t_R    g1056( .A (n1054), .Y (n1064) );
  AND2x2_ASAP7_75t_R   g1057( .A (n1064), .B (y3274), .Y (y320) );
  AO21x1_ASAP7_75t_R   g1058( .A1 (n16), .A2 (y2079), .B (x0), .Y (n1066) );
  AO21x1_ASAP7_75t_R   g1059( .A1 (n396), .A2 (n1066), .B (n581), .Y (y321) );
  OR3x1_ASAP7_75t_R    g1060( .A (n29), .B (n31), .C (n12), .Y (n1068) );
  AND2x2_ASAP7_75t_R   g1061( .A (n1068), .B (n219), .Y (y322) );
  AND2x2_ASAP7_75t_R   g1062( .A (y3274), .B (n455), .Y (y323) );
  INVx1_ASAP7_75t_R    g1063( .A (n697), .Y (n1071) );
  OR3x1_ASAP7_75t_R    g1064( .A (n1071), .B (n977), .C (n974), .Y (y324) );
  OR3x1_ASAP7_75t_R    g1065( .A (n977), .B (y2079), .C (n974), .Y (y2607) );
  AND2x2_ASAP7_75t_R   g1066( .A (y2607), .B (n445), .Y (y325) );
  NOR2x1_ASAP7_75t_R   g1067( .A (n58), .B (n466), .Y (n1075) );
  AO21x1_ASAP7_75t_R   g1068( .A1 (n466), .A2 (y2389), .B (n1075), .Y (y326) );
  AO21x1_ASAP7_75t_R   g1069( .A1 (n16), .A2 (x4), .B (x0), .Y (n1077) );
  AND2x2_ASAP7_75t_R   g1070( .A (n436), .B (y2079), .Y (n1078) );
  AO21x1_ASAP7_75t_R   g1071( .A1 (n968), .A2 (n1077), .B (n1078), .Y (y327) );
  AND2x2_ASAP7_75t_R   g1072( .A (n913), .B (x4), .Y (n1080) );
  AO21x1_ASAP7_75t_R   g1073( .A1 (n916), .A2 (x0), .B (n1080), .Y (y328) );
  AO21x1_ASAP7_75t_R   g1074( .A1 (n22), .A2 (x5), .B (x1), .Y (n1082) );
  AND2x2_ASAP7_75t_R   g1075( .A (n1082), .B (x0), .Y (n1083) );
  AO21x1_ASAP7_75t_R   g1076( .A1 (n913), .A2 (x4), .B (n1083), .Y (y329) );
  AO21x1_ASAP7_75t_R   g1077( .A1 (n466), .A2 (n58), .B (n1078), .Y (y3602) );
  AO21x1_ASAP7_75t_R   g1078( .A1 (n12), .A2 (n961), .B (y3602), .Y (y330) );
  INVx1_ASAP7_75t_R    g1079( .A (n466), .Y (n1087) );
  OA21x2_ASAP7_75t_R   g1080( .A1 (n1087), .A2 (y195), .B (n1001), .Y (y331) );
  AO21x1_ASAP7_75t_R   g1081( .A1 (n22), .A2 (x0), .B (y2079), .Y (y1281) );
  AND3x1_ASAP7_75t_R   g1082( .A (n219), .B (n90), .C (x4), .Y (n1090) );
  AO21x1_ASAP7_75t_R   g1083( .A1 (n451), .A2 (y1281), .B (n1090), .Y (y332) );
  AO21x1_ASAP7_75t_R   g1084( .A1 (y2079), .A2 (x1), .B (n12), .Y (n1092) );
  INVx1_ASAP7_75t_R    g1085( .A (n1092), .Y (n1093) );
  AO21x1_ASAP7_75t_R   g1086( .A1 (n466), .A2 (n1093), .B (n1080), .Y (y333) );
  AND3x1_ASAP7_75t_R   g1087( .A (n16), .B (y2079), .C (x4), .Y (n1095) );
  NAND2x1_ASAP7_75t_R  g1088( .A (x0), .B (n1095), .Y (n1096) );
  AND2x2_ASAP7_75t_R   g1089( .A (n1096), .B (y3852), .Y (y334) );
  AO21x1_ASAP7_75t_R   g1090( .A1 (n466), .A2 (n58), .B (n529), .Y (y633) );
  AO21x1_ASAP7_75t_R   g1091( .A1 (n43), .A2 (n28), .B (y633), .Y (y335) );
  AO21x1_ASAP7_75t_R   g1092( .A1 (n466), .A2 (n58), .B (n1080), .Y (y336) );
  OR3x1_ASAP7_75t_R    g1093( .A (n529), .B (n442), .C (x0), .Y (y337) );
  NAND2x1_ASAP7_75t_R  g1094( .A (n16), .B (n493), .Y (n1102) );
  AO21x1_ASAP7_75t_R   g1095( .A1 (x4), .A2 (n16), .B (y3852), .Y (n1103) );
  INVx1_ASAP7_75t_R    g1096( .A (n352), .Y (y2196) );
  AO21x1_ASAP7_75t_R   g1097( .A1 (n1102), .A2 (n1103), .B (y2196), .Y (y338) );
  AO21x1_ASAP7_75t_R   g1098( .A1 (n12), .A2 (n16), .B (x5), .Y (n1106) );
  NAND2x1_ASAP7_75t_R  g1099( .A (n976), .B (n1106), .Y (y2852) );
  AO21x1_ASAP7_75t_R   g1100( .A1 (x4), .A2 (n978), .B (y2852), .Y (y339) );
  AND2x2_ASAP7_75t_R   g1101( .A (n299), .B (n310), .Y (n1109) );
  INVx1_ASAP7_75t_R    g1102( .A (n1109), .Y (n1110) );
  AO21x1_ASAP7_75t_R   g1103( .A1 (n299), .A2 (n310), .B (x5), .Y (n1111) );
  OAI21x1_ASAP7_75t_R  g1104( .A1 (y2079), .A2 (n1110), .B (n1111), .Y (n1112) );
  OAI21x1_ASAP7_75t_R  g1105( .A1 (x1), .A2 (n1112), .B (n988), .Y (y340) );
  AO21x1_ASAP7_75t_R   g1106( .A1 (x0), .A2 (y2079), .B (n466), .Y (n1114) );
  NAND2x1_ASAP7_75t_R  g1107( .A (n484), .B (n439), .Y (n1115) );
  XNOR2x2_ASAP7_75t_R  g1108( .A (n1114), .B (n1115), .Y (y341) );
  NAND2x1_ASAP7_75t_R  g1109( .A (x4), .B (n781), .Y (n1117) );
  AND2x2_ASAP7_75t_R   g1110( .A (y3852), .B (n352), .Y (n1118) );
  AO32x1_ASAP7_75t_R   g1111( .A1 (n913), .A2 (x4), .A3 (n583), .B1 (n1117), .B2 (n1118), .Y (y342) );
  AO21x1_ASAP7_75t_R   g1112( .A1 (n312), .A2 (n497), .B (n22), .Y (n1120) );
  AO21x1_ASAP7_75t_R   g1113( .A1 (n16), .A2 (y2079), .B (n22), .Y (n1121) );
  INVx1_ASAP7_75t_R    g1114( .A (n1121), .Y (n1122) );
  AO32x1_ASAP7_75t_R   g1115( .A1 (x0), .A2 (n1120), .A3 (n312), .B1 (n913), .B2 (n1122), .Y (y343) );
  AND2x2_ASAP7_75t_R   g1116( .A (n1103), .B (n968), .Y (y344) );
  AO21x1_ASAP7_75t_R   g1117( .A1 (x5), .A2 (n22), .B (n90), .Y (n1125) );
  AND2x2_ASAP7_75t_R   g1118( .A (n1103), .B (n1125), .Y (y345) );
  OR3x1_ASAP7_75t_R    g1119( .A (n1090), .B (n300), .C (n495), .Y (y346) );
  INVx1_ASAP7_75t_R    g1120( .A (n1082), .Y (n1128) );
  OA21x2_ASAP7_75t_R   g1121( .A1 (n1128), .A2 (n604), .B (n968), .Y (y347) );
  OA21x2_ASAP7_75t_R   g1122( .A1 (n1128), .A2 (n604), .B (n1125), .Y (y348) );
  AO32x1_ASAP7_75t_R   g1123( .A1 (x0), .A2 (n546), .A3 (n466), .B1 (n534), .B2 (n965), .Y (y349) );
  AND2x2_ASAP7_75t_R   g1124( .A (n1000), .B (x0), .Y (n1132) );
  AO21x1_ASAP7_75t_R   g1125( .A1 (n534), .A2 (n965), .B (n1132), .Y (y350) );
  NOR2x1_ASAP7_75t_R   g1126( .A (n43), .B (n137), .Y (n1134) );
  AO21x1_ASAP7_75t_R   g1127( .A1 (n56), .A2 (x3), .B (n1134), .Y (n1135) );
  NAND2x1_ASAP7_75t_R  g1128( .A (n144), .B (n1135), .Y (y351) );
  AND3x1_ASAP7_75t_R   g1129( .A (x0), .B (x4), .C (x5), .Y (n1137) );
  INVx1_ASAP7_75t_R    g1130( .A (n1137), .Y (n1138) );
  INVx1_ASAP7_75t_R    g1131( .A (n565), .Y (n1139) );
  AND3x1_ASAP7_75t_R   g1132( .A (n455), .B (y3852), .C (x1), .Y (n1140) );
  AO21x1_ASAP7_75t_R   g1133( .A1 (n1138), .A2 (n1139), .B (n1140), .Y (y352) );
  AND2x2_ASAP7_75t_R   g1134( .A (n466), .B (y3852), .Y (y3127) );
  AO21x1_ASAP7_75t_R   g1135( .A1 (y3127), .A2 (n546), .B (n974), .Y (y353) );
  OR3x1_ASAP7_75t_R    g1136( .A (n45), .B (x0), .C (x1), .Y (n1144) );
  INVx1_ASAP7_75t_R    g1137( .A (n1144), .Y (n1145) );
  NOR2x1_ASAP7_75t_R   g1138( .A (n125), .B (n63), .Y (n1146) );
  NOR2x1_ASAP7_75t_R   g1139( .A (n1145), .B (n1146), .Y (y354) );
  AND2x2_ASAP7_75t_R   g1140( .A (n1000), .B (y3852), .Y (y1775) );
  AO21x1_ASAP7_75t_R   g1141( .A1 (n28), .A2 (n43), .B (y1775), .Y (y355) );
  AND3x1_ASAP7_75t_R   g1142( .A (n22), .B (x1), .C (x0), .Y (n1150) );
  INVx1_ASAP7_75t_R    g1143( .A (n1150), .Y (n1151) );
  AO32x1_ASAP7_75t_R   g1144( .A1 (y2079), .A2 (n1151), .A3 (n466), .B1 (n299), .B2 (n594), .Y (y356) );
  AND3x1_ASAP7_75t_R   g1145( .A (n1103), .B (n968), .C (n455), .Y (y357) );
  NAND2x1_ASAP7_75t_R  g1146( .A (x4), .B (n978), .Y (n1154) );
  INVx1_ASAP7_75t_R    g1147( .A (n1154), .Y (n1155) );
  OR3x1_ASAP7_75t_R    g1148( .A (n1155), .B (n977), .C (n495), .Y (y358) );
  AND2x2_ASAP7_75t_R   g1149( .A (n1102), .B (n917), .Y (y359) );
  INVx1_ASAP7_75t_R    g1150( .A (n360), .Y (n1158) );
  OR3x1_ASAP7_75t_R    g1151( .A (n1158), .B (n291), .C (y3852), .Y (y1308) );
  AND3x1_ASAP7_75t_R   g1152( .A (n671), .B (n22), .C (x0), .Y (n1160) );
  INVx1_ASAP7_75t_R    g1153( .A (n1160), .Y (n1161) );
  AND2x2_ASAP7_75t_R   g1154( .A (y1308), .B (n1161), .Y (y360) );
  AO21x1_ASAP7_75t_R   g1155( .A1 (y2079), .A2 (x0), .B (x4), .Y (n1163) );
  INVx1_ASAP7_75t_R    g1156( .A (n1163), .Y (n1164) );
  OA22x2_ASAP7_75t_R   g1157( .A1 (n1164), .A2 (n488), .B1 (n1128), .B2 (n604), .Y (y361) );
  AO21x1_ASAP7_75t_R   g1158( .A1 (n22), .A2 (x0), .B (x1), .Y (n1166) );
  AO21x1_ASAP7_75t_R   g1159( .A1 (n455), .A2 (x0), .B (n541), .Y (n1167) );
  OA21x2_ASAP7_75t_R   g1160( .A1 (n386), .A2 (n1166), .B (n1167), .Y (y362) );
  INVx1_ASAP7_75t_R    g1161( .A (n916), .Y (n1169) );
  OA21x2_ASAP7_75t_R   g1162( .A1 (n1169), .A2 (n1093), .B (n1102), .Y (y363) );
  AND3x1_ASAP7_75t_R   g1163( .A (n1102), .B (n1103), .C (n455), .Y (y364) );
  NAND2x1_ASAP7_75t_R  g1164( .A (n12), .B (n561), .Y (y365) );
  INVx1_ASAP7_75t_R    g1165( .A (n1000), .Y (n1173) );
  OA21x2_ASAP7_75t_R   g1166( .A1 (x0), .A2 (n1173), .B (n919), .Y (y366) );
  AO21x1_ASAP7_75t_R   g1167( .A1 (n22), .A2 (x1), .B (x0), .Y (n1175) );
  AO21x1_ASAP7_75t_R   g1168( .A1 (n466), .A2 (x0), .B (n974), .Y (n1176) );
  AO21x1_ASAP7_75t_R   g1169( .A1 (y2079), .A2 (n1175), .B (n1176), .Y (y367) );
  AND2x2_ASAP7_75t_R   g1170( .A (n919), .B (n1077), .Y (y368) );
  AO21x1_ASAP7_75t_R   g1171( .A1 (n765), .A2 (n1087), .B (n1083), .Y (y369) );
  AND3x1_ASAP7_75t_R   g1172( .A (n455), .B (n90), .C (n219), .Y (n1180) );
  AO21x1_ASAP7_75t_R   g1173( .A1 (n556), .A2 (n173), .B (n1180), .Y (y370) );
  INVx1_ASAP7_75t_R    g1174( .A (n938), .Y (n1182) );
  AO32x1_ASAP7_75t_R   g1175( .A1 (x0), .A2 (n1114), .A3 (n546), .B1 (n584), .B2 (n1182), .Y (y371) );
  AND2x2_ASAP7_75t_R   g1176( .A (n466), .B (n58), .Y (n1184) );
  AO21x1_ASAP7_75t_R   g1177( .A1 (n913), .A2 (n310), .B (n1184), .Y (y372) );
  AO21x1_ASAP7_75t_R   g1178( .A1 (n12), .A2 (x4), .B (y2079), .Y (n1186) );
  AO21x1_ASAP7_75t_R   g1179( .A1 (n16), .A2 (n1186), .B (n1132), .Y (y373) );
  AO21x1_ASAP7_75t_R   g1180( .A1 (n16), .A2 (n22), .B (x0), .Y (n1188) );
  INVx1_ASAP7_75t_R    g1181( .A (n1188), .Y (n1189) );
  AND3x1_ASAP7_75t_R   g1182( .A (n16), .B (x4), .C (x5), .Y (n1190) );
  INVx1_ASAP7_75t_R    g1183( .A (n1190), .Y (n1191) );
  AO32x1_ASAP7_75t_R   g1184( .A1 (n388), .A2 (n1189), .A3 (n776), .B1 (x0), .B2 (n1191), .Y (y374) );
  AND3x1_ASAP7_75t_R   g1185( .A (n28), .B (n388), .C (n16), .Y (n1193) );
  OAI21x1_ASAP7_75t_R  g1186( .A1 (n1193), .A2 (n12), .B (y4), .Y (y375) );
  AND3x1_ASAP7_75t_R   g1187( .A (n16), .B (x5), .C (x4), .Y (n1195) );
  INVx1_ASAP7_75t_R    g1188( .A (n1195), .Y (n1196) );
  NOR2x1_ASAP7_75t_R   g1189( .A (n1082), .B (n604), .Y (n1197) );
  AO21x1_ASAP7_75t_R   g1190( .A1 (n1196), .A2 (x0), .B (n1197), .Y (y376) );
  NOR2x1_ASAP7_75t_R   g1191( .A (n12), .B (n1195), .Y (y2778) );
  AO21x1_ASAP7_75t_R   g1192( .A1 (x5), .A2 (n974), .B (y2778), .Y (y377) );
  OR3x1_ASAP7_75t_R    g1193( .A (n29), .B (n25), .C (n12), .Y (n1201) );
  OA21x2_ASAP7_75t_R   g1194( .A1 (x0), .A2 (n1195), .B (n1201), .Y (y378) );
  AND3x1_ASAP7_75t_R   g1195( .A (n90), .B (n22), .C (y2079), .Y (n1203) );
  INVx1_ASAP7_75t_R    g1196( .A (n1203), .Y (n1204) );
  AND2x2_ASAP7_75t_R   g1197( .A (n90), .B (n22), .Y (n1205) );
  AO21x1_ASAP7_75t_R   g1198( .A1 (n1205), .A2 (y2079), .B (n1195), .Y (n1206) );
  AO32x1_ASAP7_75t_R   g1199( .A1 (n1196), .A2 (n1204), .A3 (x0), .B1 (n12), .B2 (n1206), .Y (y379) );
  INVx1_ASAP7_75t_R    g1200( .A (n219), .Y (n1208) );
  AO21x1_ASAP7_75t_R   g1201( .A1 (n16), .A2 (x0), .B (y2079), .Y (n1209) );
  INVx1_ASAP7_75t_R    g1202( .A (n1209), .Y (n1210) );
  OR3x1_ASAP7_75t_R    g1203( .A (n1208), .B (n1210), .C (x4), .Y (n1211) );
  AND2x2_ASAP7_75t_R   g1204( .A (n1211), .B (n387), .Y (y380) );
  AO21x1_ASAP7_75t_R   g1205( .A1 (n22), .A2 (n312), .B (n31), .Y (n1213) );
  INVx1_ASAP7_75t_R    g1206( .A (n1213), .Y (n1214) );
  AO21x1_ASAP7_75t_R   g1207( .A1 (y2079), .A2 (x4), .B (n544), .Y (n1215) );
  OR3x1_ASAP7_75t_R    g1208( .A (n1215), .B (n12), .C (n527), .Y (n1216) );
  OA21x2_ASAP7_75t_R   g1209( .A1 (n1214), .A2 (x0), .B (n1216), .Y (y381) );
  OR3x1_ASAP7_75t_R    g1210( .A (n544), .B (n12), .C (x4), .Y (n1218) );
  AND2x2_ASAP7_75t_R   g1211( .A (n387), .B (n1218), .Y (y382) );
  AO21x1_ASAP7_75t_R   g1212( .A1 (n28), .A2 (n30), .B (x0), .Y (n1220) );
  AND2x2_ASAP7_75t_R   g1213( .A (n1068), .B (n1220), .Y (y383) );
  NAND2x1_ASAP7_75t_R  g1214( .A (n16), .B (n430), .Y (n1222) );
  INVx1_ASAP7_75t_R    g1215( .A (n1222), .Y (n1223) );
  AO21x1_ASAP7_75t_R   g1216( .A1 (n613), .A2 (n1223), .B (y689), .Y (y384) );
  OA21x2_ASAP7_75t_R   g1217( .A1 (x0), .A2 (n1193), .B (n1068), .Y (y385) );
  AND3x1_ASAP7_75t_R   g1218( .A (n90), .B (n219), .C (x5), .Y (n1226) );
  AO21x1_ASAP7_75t_R   g1219( .A1 (y2079), .A2 (n175), .B (n1226), .Y (y386) );
  AO21x1_ASAP7_75t_R   g1220( .A1 (y2079), .A2 (y25), .B (y232), .Y (y387) );
  AO21x1_ASAP7_75t_R   g1221( .A1 (y2079), .A2 (x2), .B (n143), .Y (n1229) );
  AO21x1_ASAP7_75t_R   g1222( .A1 (n481), .A2 (n16), .B (n1229), .Y (y388) );
  AND3x1_ASAP7_75t_R   g1223( .A (n15), .B (x0), .C (x1), .Y (n1231) );
  INVx1_ASAP7_75t_R    g1224( .A (n1231), .Y (n1232) );
  AO21x1_ASAP7_75t_R   g1225( .A1 (y2079), .A2 (n1232), .B (n1226), .Y (y389) );
  AND3x1_ASAP7_75t_R   g1226( .A (n90), .B (n219), .C (n15), .Y (n1234) );
  NAND2x1_ASAP7_75t_R  g1227( .A (y2079), .B (n1234), .Y (n1235) );
  AND2x2_ASAP7_75t_R   g1228( .A (n1235), .B (y1873), .Y (y390) );
  AND3x1_ASAP7_75t_R   g1229( .A (n90), .B (y2079), .C (n15), .Y (n1237) );
  INVx1_ASAP7_75t_R    g1230( .A (n908), .Y (n1238) );
  NOR2x1_ASAP7_75t_R   g1231( .A (n1237), .B (n1238), .Y (y391) );
  INVx1_ASAP7_75t_R    g1232( .A (n950), .Y (n1240) );
  AO21x1_ASAP7_75t_R   g1233( .A1 (y2079), .A2 (n1240), .B (n1226), .Y (y392) );
  AO21x1_ASAP7_75t_R   g1234( .A1 (n16), .A2 (n12), .B (x5), .Y (n1242) );
  INVx1_ASAP7_75t_R    g1235( .A (n1242), .Y (y2093) );
  OR3x1_ASAP7_75t_R    g1236( .A (y2093), .B (n38), .C (y863), .Y (y393) );
  AND3x1_ASAP7_75t_R   g1237( .A (n16), .B (x5), .C (x0), .Y (n1245) );
  INVx1_ASAP7_75t_R    g1238( .A (n1245), .Y (n1246) );
  AO21x1_ASAP7_75t_R   g1239( .A1 (n16), .A2 (x5), .B (x0), .Y (n1247) );
  AND3x1_ASAP7_75t_R   g1240( .A (y2079), .B (x2), .C (x1), .Y (n1248) );
  AO21x1_ASAP7_75t_R   g1241( .A1 (n1246), .A2 (n1247), .B (n1248), .Y (y394) );
  AO21x1_ASAP7_75t_R   g1242( .A1 (y9), .A2 (n746), .B (n128), .Y (n1250) );
  NOR2x1_ASAP7_75t_R   g1243( .A (x5), .B (n1250), .Y (n1251) );
  NOR2x1_ASAP7_75t_R   g1244( .A (n1238), .B (n1251), .Y (y395) );
  AND3x1_ASAP7_75t_R   g1245( .A (n12), .B (n16), .C (x3), .Y (n1253) );
  AO21x1_ASAP7_75t_R   g1246( .A1 (n12), .A2 (x3), .B (n16), .Y (n1254) );
  INVx1_ASAP7_75t_R    g1247( .A (n1254), .Y (n1255) );
  OA33x2_ASAP7_75t_R   g1248( .A1 (n15), .A2 (n243), .A3 (x0), .B1 (x2), .B2 (n1253), .B3 (n1255), .Y (y396) );
  AO21x1_ASAP7_75t_R   g1249( .A1 (n15), .A2 (x0), .B (n16), .Y (n1257) );
  AND3x1_ASAP7_75t_R   g1250( .A (n90), .B (n1257), .C (y2079), .Y (n1258) );
  INVx1_ASAP7_75t_R    g1251( .A (y1873), .Y (n1259) );
  NOR2x1_ASAP7_75t_R   g1252( .A (n1258), .B (n1259), .Y (y397) );
  INVx1_ASAP7_75t_R    g1253( .A (n63), .Y (n1261) );
  INVx1_ASAP7_75t_R    g1254( .A (n64), .Y (n1262) );
  OR3x1_ASAP7_75t_R    g1255( .A (n1261), .B (n1262), .C (n84), .Y (n1263) );
  NAND2x1_ASAP7_75t_R  g1256( .A (n155), .B (n1263), .Y (y398) );
  INVx1_ASAP7_75t_R    g1257( .A (n856), .Y (n1265) );
  AND3x1_ASAP7_75t_R   g1258( .A (n1265), .B (y3852), .C (x1), .Y (n1266) );
  AO21x1_ASAP7_75t_R   g1259( .A1 (n765), .A2 (n1139), .B (n1266), .Y (y399) );
  AO21x1_ASAP7_75t_R   g1260( .A1 (n348), .A2 (x0), .B (y2723), .Y (y400) );
  INVx1_ASAP7_75t_R    g1261( .A (n740), .Y (n1269) );
  AO21x1_ASAP7_75t_R   g1262( .A1 (n228), .A2 (n1269), .B (n1226), .Y (y401) );
  NAND2x1_ASAP7_75t_R  g1263( .A (x0), .B (n1050), .Y (n1271) );
  OR3x1_ASAP7_75t_R    g1264( .A (y2466), .B (n16), .C (x0), .Y (n1272) );
  AO21x1_ASAP7_75t_R   g1265( .A1 (n1271), .A2 (n1272), .B (y2196), .Y (y402) );
  AND2x2_ASAP7_75t_R   g1266( .A (n445), .B (n1047), .Y (y403) );
  AO21x1_ASAP7_75t_R   g1267( .A1 (x4), .A2 (y2079), .B (n90), .Y (n1275) );
  AND2x2_ASAP7_75t_R   g1268( .A (n1275), .B (n1272), .Y (y404) );
  AND3x1_ASAP7_75t_R   g1269( .A (n17), .B (x4), .C (x5), .Y (n1277) );
  AO21x1_ASAP7_75t_R   g1270( .A1 (n22), .A2 (n319), .B (n1277), .Y (n1278) );
  OR3x1_ASAP7_75t_R    g1271( .A (n1278), .B (n537), .C (n628), .Y (y405) );
  NAND2x1_ASAP7_75t_R  g1272( .A (n1103), .B (n1102), .Y (n1280) );
  INVx1_ASAP7_75t_R    g1273( .A (n1280), .Y (y3445) );
  OR3x1_ASAP7_75t_R    g1274( .A (y3445), .B (y2196), .C (n437), .Y (y406) );
  AO21x1_ASAP7_75t_R   g1275( .A1 (n455), .A2 (n765), .B (x1), .Y (n1283) );
  AND2x2_ASAP7_75t_R   g1276( .A (n1283), .B (n1272), .Y (y407) );
  NOR2x1_ASAP7_75t_R   g1277( .A (n1245), .B (n1208), .Y (y408) );
  AO21x1_ASAP7_75t_R   g1278( .A1 (n1265), .A2 (n43), .B (y772), .Y (y409) );
  AO21x1_ASAP7_75t_R   g1279( .A1 (n1265), .A2 (n765), .B (x1), .Y (n1287) );
  AND2x2_ASAP7_75t_R   g1280( .A (n1287), .B (n219), .Y (y410) );
  OR3x1_ASAP7_75t_R    g1281( .A (n143), .B (x5), .C (x2), .Y (n1289) );
  INVx1_ASAP7_75t_R    g1282( .A (n1289), .Y (n1290) );
  OR3x1_ASAP7_75t_R    g1283( .A (n856), .B (n16), .C (n12), .Y (n1291) );
  INVx1_ASAP7_75t_R    g1284( .A (n1291), .Y (n1292) );
  OR3x1_ASAP7_75t_R    g1285( .A (n1290), .B (n1060), .C (n1292), .Y (y411) );
  AO21x1_ASAP7_75t_R   g1286( .A1 (n84), .A2 (x1), .B (n1253), .Y (n1294) );
  NAND2x1_ASAP7_75t_R  g1287( .A (x1), .B (n17), .Y (n1295) );
  NAND2x1_ASAP7_75t_R  g1288( .A (x3), .B (n16), .Y (n1296) );
  AND2x2_ASAP7_75t_R   g1289( .A (n1295), .B (n1296), .Y (n1297) );
  OA22x2_ASAP7_75t_R   g1290( .A1 (x2), .A2 (n1294), .B1 (n1297), .B2 (n244), .Y (y412) );
  AND2x2_ASAP7_75t_R   g1291( .A (n219), .B (n90), .Y (n1299) );
  INVx1_ASAP7_75t_R    g1292( .A (n1299), .Y (n1300) );
  AO21x1_ASAP7_75t_R   g1293( .A1 (n16), .A2 (x0), .B (n15), .Y (n1301) );
  AND2x2_ASAP7_75t_R   g1294( .A (n1301), .B (y2079), .Y (n1302) );
  AND3x1_ASAP7_75t_R   g1295( .A (n1265), .B (n219), .C (n90), .Y (n1303) );
  AO21x1_ASAP7_75t_R   g1296( .A1 (n1300), .A2 (n1302), .B (n1303), .Y (y413) );
  AO21x1_ASAP7_75t_R   g1297( .A1 (n16), .A2 (n12), .B (y2079), .Y (n1305) );
  INVx1_ASAP7_75t_R    g1298( .A (n905), .Y (n1306) );
  AO32x1_ASAP7_75t_R   g1299( .A1 (n466), .A2 (n1175), .A3 (x5), .B1 (n1305), .B2 (n1306), .Y (y414) );
  AND2x2_ASAP7_75t_R   g1300( .A (n665), .B (x0), .Y (y890) );
  AO21x1_ASAP7_75t_R   g1301( .A1 (n12), .A2 (n758), .B (y890), .Y (y415) );
  NAND2x1_ASAP7_75t_R  g1302( .A (n22), .B (n1305), .Y (n1310) );
  AO21x1_ASAP7_75t_R   g1303( .A1 (x1), .A2 (x0), .B (x5), .Y (n1311) );
  INVx1_ASAP7_75t_R    g1304( .A (n1311), .Y (n1312) );
  AO21x1_ASAP7_75t_R   g1305( .A1 (n899), .A2 (n1310), .B (n1312), .Y (y416) );
  AND2x2_ASAP7_75t_R   g1306( .A (n1265), .B (n219), .Y (n1314) );
  AND3x1_ASAP7_75t_R   g1307( .A (n241), .B (y2079), .C (x1), .Y (n1315) );
  AO21x1_ASAP7_75t_R   g1308( .A1 (n1314), .A2 (n1246), .B (n1315), .Y (y417) );
  AND3x1_ASAP7_75t_R   g1309( .A (x2), .B (x1), .C (x3), .Y (n1317) );
  OR3x1_ASAP7_75t_R    g1310( .A (y1081), .B (n1317), .C (n109), .Y (y418) );
  AO21x1_ASAP7_75t_R   g1311( .A1 (x0), .A2 (x3), .B (x4), .Y (n1319) );
  AND2x2_ASAP7_75t_R   g1312( .A (n624), .B (n1319), .Y (n1320) );
  AO21x1_ASAP7_75t_R   g1313( .A1 (n352), .A2 (n337), .B (n1320), .Y (y419) );
  AO21x1_ASAP7_75t_R   g1314( .A1 (y2079), .A2 (x2), .B (n43), .Y (n1322) );
  AO21x1_ASAP7_75t_R   g1315( .A1 (x1), .A2 (n58), .B (n1322), .Y (y3940) );
  NAND2x1_ASAP7_75t_R  g1316( .A (n12), .B (n705), .Y (n1324) );
  AND2x2_ASAP7_75t_R   g1317( .A (y3940), .B (n1324), .Y (y420) );
  AO21x1_ASAP7_75t_R   g1318( .A1 (n776), .A2 (n388), .B (x0), .Y (n1326) );
  AND2x2_ASAP7_75t_R   g1319( .A (n1326), .B (n1246), .Y (y421) );
  AND3x1_ASAP7_75t_R   g1320( .A (y103), .B (n505), .C (n419), .Y (y422) );
  AND3x1_ASAP7_75t_R   g1321( .A (n388), .B (n219), .C (n90), .Y (n1329) );
  AO21x1_ASAP7_75t_R   g1322( .A1 (y2079), .A2 (x0), .B (n1329), .Y (y423) );
  OR3x1_ASAP7_75t_R    g1323( .A (n1269), .B (n12), .C (n544), .Y (n1331) );
  AO21x1_ASAP7_75t_R   g1324( .A1 (n776), .A2 (n740), .B (x0), .Y (n1332) );
  AND2x2_ASAP7_75t_R   g1325( .A (n1331), .B (n1332), .Y (y424) );
  AO21x1_ASAP7_75t_R   g1326( .A1 (n388), .A2 (n28), .B (n125), .Y (n1334) );
  OA21x2_ASAP7_75t_R   g1327( .A1 (y3758), .A2 (n84), .B (n1334), .Y (y425) );
  AO21x1_ASAP7_75t_R   g1328( .A1 (y2079), .A2 (x2), .B (x1), .Y (n1336) );
  INVx1_ASAP7_75t_R    g1329( .A (n1336), .Y (n1337) );
  AO21x1_ASAP7_75t_R   g1330( .A1 (n692), .A2 (n1337), .B (y890), .Y (y426) );
  AND3x1_ASAP7_75t_R   g1331( .A (n15), .B (y2079), .C (x1), .Y (n1339) );
  INVx1_ASAP7_75t_R    g1332( .A (n1339), .Y (n1340) );
  AND3x1_ASAP7_75t_R   g1333( .A (n1340), .B (n1246), .C (n1247), .Y (y427) );
  AO21x1_ASAP7_75t_R   g1334( .A1 (x3), .A2 (x4), .B (x0), .Y (n1342) );
  INVx1_ASAP7_75t_R    g1335( .A (n1342), .Y (n1343) );
  AO21x1_ASAP7_75t_R   g1336( .A1 (n639), .A2 (n1343), .B (n1320), .Y (y428) );
  AO21x1_ASAP7_75t_R   g1337( .A1 (n740), .A2 (n16), .B (x0), .Y (n1345) );
  AND2x2_ASAP7_75t_R   g1338( .A (n1331), .B (n1345), .Y (y429) );
  AO21x1_ASAP7_75t_R   g1339( .A1 (n665), .A2 (x0), .B (n978), .Y (y430) );
  AO21x1_ASAP7_75t_R   g1340( .A1 (n90), .A2 (n219), .B (y2466), .Y (y431) );
  INVx1_ASAP7_75t_R    g1341( .A (y8), .Y (n1349) );
  INVx1_ASAP7_75t_R    g1342( .A (n453), .Y (y2482) );
  OR3x1_ASAP7_75t_R    g1343( .A (n1349), .B (y2482), .C (n143), .Y (y432) );
  INVx1_ASAP7_75t_R    g1344( .A (n781), .Y (n1352) );
  AO21x1_ASAP7_75t_R   g1345( .A1 (n1352), .A2 (n22), .B (n493), .Y (y433) );
  OR3x1_ASAP7_75t_R    g1346( .A (n315), .B (x5), .C (x1), .Y (n1354) );
  AND2x2_ASAP7_75t_R   g1347( .A (n1354), .B (y3852), .Y (y434) );
  OR3x1_ASAP7_75t_R    g1348( .A (y863), .B (x3), .C (x2), .Y (n1356) );
  INVx1_ASAP7_75t_R    g1349( .A (n1356), .Y (n1357) );
  OR3x1_ASAP7_75t_R    g1350( .A (n45), .B (n12), .C (n16), .Y (n1358) );
  INVx1_ASAP7_75t_R    g1351( .A (n1358), .Y (n1359) );
  OR3x1_ASAP7_75t_R    g1352( .A (n1357), .B (n1359), .C (n227), .Y (y436) );
  AND3x1_ASAP7_75t_R   g1353( .A (n168), .B (n167), .C (n16), .Y (n1361) );
  INVx1_ASAP7_75t_R    g1354( .A (n168), .Y (n1362) );
  INVx1_ASAP7_75t_R    g1355( .A (n167), .Y (n1363) );
  OA21x2_ASAP7_75t_R   g1356( .A1 (n1362), .A2 (n1363), .B (x1), .Y (n1364) );
  OR2x4_ASAP7_75t_R    g1357( .A (n1361), .B (n1364), .Y (y437) );
  AO21x1_ASAP7_75t_R   g1358( .A1 (n1062), .A2 (n143), .B (n43), .Y (y438) );
  AND3x1_ASAP7_75t_R   g1359( .A (n1062), .B (n90), .C (n219), .Y (y439) );
  OR3x1_ASAP7_75t_R    g1360( .A (n186), .B (y2079), .C (y863), .Y (y440) );
  AND3x1_ASAP7_75t_R   g1361( .A (y2079), .B (n22), .C (x0), .Y (y2498) );
  INVx1_ASAP7_75t_R    g1362( .A (y2498), .Y (n1370) );
  AND2x2_ASAP7_75t_R   g1363( .A (y116), .B (n1370), .Y (y441) );
  AO21x1_ASAP7_75t_R   g1364( .A1 (n1305), .A2 (n175), .B (y863), .Y (y442) );
  AO21x1_ASAP7_75t_R   g1365( .A1 (n12), .A2 (x2), .B (y2079), .Y (n1373) );
  AO22x1_ASAP7_75t_R   g1366( .A1 (n16), .A2 (n1373), .B1 (x1), .B2 (n707), .Y (y443) );
  AO21x1_ASAP7_75t_R   g1367( .A1 (n1305), .A2 (x2), .B (y863), .Y (y444) );
  AND3x1_ASAP7_75t_R   g1368( .A (n90), .B (n219), .C (n800), .Y (n1376) );
  AO21x1_ASAP7_75t_R   g1369( .A1 (n221), .A2 (y2079), .B (n1376), .Y (y445) );
  AO21x1_ASAP7_75t_R   g1370( .A1 (y9), .A2 (n312), .B (x2), .Y (n1378) );
  AND2x2_ASAP7_75t_R   g1371( .A (n1378), .B (n908), .Y (y446) );
  AND3x1_ASAP7_75t_R   g1372( .A (x1), .B (x0), .C (x5), .Y (n1380) );
  AO21x1_ASAP7_75t_R   g1373( .A1 (y2079), .A2 (x2), .B (n1380), .Y (y2155) );
  AO21x1_ASAP7_75t_R   g1374( .A1 (n227), .A2 (n97), .B (y2155), .Y (y447) );
  AO21x1_ASAP7_75t_R   g1375( .A1 (y2079), .A2 (n244), .B (n989), .Y (n1383) );
  AO21x1_ASAP7_75t_R   g1376( .A1 (x2), .A2 (n978), .B (n1383), .Y (y448) );
  OR3x1_ASAP7_75t_R    g1377( .A (x1), .B (x0), .C (x5), .Y (n1385) );
  AND2x2_ASAP7_75t_R   g1378( .A (y440), .B (n1385), .Y (y449) );
  INVx1_ASAP7_75t_R    g1379( .A (n701), .Y (n1387) );
  AO32x1_ASAP7_75t_R   g1380( .A1 (n16), .A2 (n1373), .A3 (n1387), .B1 (x1), .B2 (n707), .Y (y450) );
  AO21x1_ASAP7_75t_R   g1381( .A1 (n312), .A2 (n497), .B (n15), .Y (n1389) );
  AOI21x1_ASAP7_75t_R  g1382( .A1 (n12), .A2 (n1389), .B (n1245), .Y (y451) );
  AO21x1_ASAP7_75t_R   g1383( .A1 (n16), .A2 (n12), .B (x2), .Y (n1391) );
  AO21x1_ASAP7_75t_R   g1384( .A1 (n1391), .A2 (y2079), .B (y863), .Y (y1283) );
  NAND2x1_ASAP7_75t_R  g1385( .A (n16), .B (n701), .Y (n1393) );
  OA21x2_ASAP7_75t_R   g1386( .A1 (n186), .A2 (y1283), .B (n1393), .Y (y452) );
  AND2x2_ASAP7_75t_R   g1387( .A (y444), .B (n1385), .Y (y453) );
  OR3x1_ASAP7_75t_R    g1388( .A (n291), .B (n293), .C (x0), .Y (y454) );
  AO21x1_ASAP7_75t_R   g1389( .A1 (x1), .A2 (x0), .B (n186), .Y (y2393) );
  AO32x1_ASAP7_75t_R   g1390( .A1 (y2079), .A2 (n1232), .A3 (n228), .B1 (x5), .B2 (y2393), .Y (y455) );
  AND3x1_ASAP7_75t_R   g1391( .A (x0), .B (x5), .C (x4), .Y (n1399) );
  INVx1_ASAP7_75t_R    g1392( .A (n1399), .Y (n1400) );
  AO32x1_ASAP7_75t_R   g1393( .A1 (n16), .A2 (n419), .A3 (n1400), .B1 (x1), .B2 (y1894), .Y (y456) );
  INVx1_ASAP7_75t_R    g1394( .A (n747), .Y (n1402) );
  AO21x1_ASAP7_75t_R   g1395( .A1 (x1), .A2 (x2), .B (x5), .Y (n1403) );
  AND3x1_ASAP7_75t_R   g1396( .A (n12), .B (n16), .C (x2), .Y (n1404) );
  OR3x1_ASAP7_75t_R    g1397( .A (n1404), .B (y2079), .C (n143), .Y (n1405) );
  OA21x2_ASAP7_75t_R   g1398( .A1 (n1402), .A2 (n1403), .B (n1405), .Y (y457) );
  AO21x1_ASAP7_75t_R   g1399( .A1 (x1), .A2 (x5), .B (n15), .Y (n1407) );
  INVx1_ASAP7_75t_R    g1400( .A (n1407), .Y (n1408) );
  AND3x1_ASAP7_75t_R   g1401( .A (y3852), .B (n352), .C (n16), .Y (n1409) );
  INVx1_ASAP7_75t_R    g1402( .A (n1409), .Y (n1410) );
  OA21x2_ASAP7_75t_R   g1403( .A1 (n1408), .A2 (n1093), .B (n1410), .Y (y458) );
  AND3x1_ASAP7_75t_R   g1404( .A (n187), .B (n1391), .C (y2079), .Y (n1412) );
  AO21x1_ASAP7_75t_R   g1405( .A1 (y2393), .A2 (x5), .B (n1412), .Y (y459) );
  NOR2x1_ASAP7_75t_R   g1406( .A (n227), .B (n740), .Y (n1414) );
  AO21x1_ASAP7_75t_R   g1407( .A1 (y2393), .A2 (x5), .B (n1414), .Y (y460) );
  AO21x1_ASAP7_75t_R   g1408( .A1 (n15), .A2 (y2079), .B (n143), .Y (n1416) );
  AO21x1_ASAP7_75t_R   g1409( .A1 (n1262), .A2 (n765), .B (n1416), .Y (y461) );
  AO21x1_ASAP7_75t_R   g1410( .A1 (n994), .A2 (n858), .B (n1404), .Y (y462) );
  NOR2x1_ASAP7_75t_R   g1411( .A (n58), .B (n64), .Y (n1419) );
  AO21x1_ASAP7_75t_R   g1412( .A1 (n858), .A2 (x1), .B (n1419), .Y (y463) );
  NOR2x1_ASAP7_75t_R   g1413( .A (x0), .B (n602), .Y (n1421) );
  INVx1_ASAP7_75t_R    g1414( .A (n1421), .Y (n1422) );
  AND2x2_ASAP7_75t_R   g1415( .A (n1422), .B (y370), .Y (y464) );
  AO21x1_ASAP7_75t_R   g1416( .A1 (n16), .A2 (x2), .B (x0), .Y (n1424) );
  AND2x2_ASAP7_75t_R   g1417( .A (n1246), .B (n1424), .Y (y465) );
  AO21x1_ASAP7_75t_R   g1418( .A1 (n12), .A2 (n15), .B (n16), .Y (n1426) );
  AO21x1_ASAP7_75t_R   g1419( .A1 (n1426), .A2 (n1373), .B (n1292), .Y (y466) );
  AO21x1_ASAP7_75t_R   g1420( .A1 (n15), .A2 (x5), .B (n103), .Y (n1428) );
  INVx1_ASAP7_75t_R    g1421( .A (n1428), .Y (n1429) );
  AO21x1_ASAP7_75t_R   g1422( .A1 (n12), .A2 (n1429), .B (y890), .Y (y467) );
  AO21x1_ASAP7_75t_R   g1423( .A1 (n12), .A2 (y2079), .B (x3), .Y (n1431) );
  INVx1_ASAP7_75t_R    g1424( .A (n1431), .Y (n1432) );
  OR3x1_ASAP7_75t_R    g1425( .A (n1432), .B (n299), .C (n425), .Y (n1433) );
  INVx1_ASAP7_75t_R    g1426( .A (n425), .Y (n1434) );
  AO21x1_ASAP7_75t_R   g1427( .A1 (n1434), .A2 (n1431), .B (x4), .Y (n1435) );
  AND2x2_ASAP7_75t_R   g1428( .A (n1433), .B (n1435), .Y (y468) );
  NOR2x1_ASAP7_75t_R   g1429( .A (n15), .B (n58), .Y (n1437) );
  OR3x1_ASAP7_75t_R    g1430( .A (n856), .B (n16), .C (x0), .Y (n1438) );
  OA21x2_ASAP7_75t_R   g1431( .A1 (n1437), .A2 (n1352), .B (n1438), .Y (y469) );
  AO21x1_ASAP7_75t_R   g1432( .A1 (x2), .A2 (n12), .B (n497), .Y (n1440) );
  AND3x1_ASAP7_75t_R   g1433( .A (n1440), .B (n714), .C (n219), .Y (y470) );
  AND2x2_ASAP7_75t_R   g1434( .A (y630), .B (n455), .Y (y471) );
  AND2x2_ASAP7_75t_R   g1435( .A (n1247), .B (n747), .Y (n1443) );
  AO21x1_ASAP7_75t_R   g1436( .A1 (y2079), .A2 (n244), .B (n1443), .Y (y472) );
  AND2x2_ASAP7_75t_R   g1437( .A (n858), .B (n994), .Y (n1445) );
  AO21x1_ASAP7_75t_R   g1438( .A1 (x2), .A2 (n978), .B (n1445), .Y (y473) );
  OA21x2_ASAP7_75t_R   g1439( .A1 (n128), .A2 (n1247), .B (n1440), .Y (y474) );
  AND2x2_ASAP7_75t_R   g1440( .A (n844), .B (y3852), .Y (y475) );
  OA21x2_ASAP7_75t_R   g1441( .A1 (n1437), .A2 (x1), .B (n1345), .Y (y476) );
  AO21x1_ASAP7_75t_R   g1442( .A1 (n16), .A2 (x2), .B (y2079), .Y (n1450) );
  AO21x1_ASAP7_75t_R   g1443( .A1 (n740), .A2 (n1450), .B (x0), .Y (n1451) );
  AND2x2_ASAP7_75t_R   g1444( .A (n1331), .B (n1451), .Y (y477) );
  AO21x1_ASAP7_75t_R   g1445( .A1 (x0), .A2 (x1), .B (x2), .Y (n1453) );
  INVx1_ASAP7_75t_R    g1446( .A (n1453), .Y (n1454) );
  NAND2x1_ASAP7_75t_R  g1447( .A (x5), .B (n797), .Y (n1455) );
  OA21x2_ASAP7_75t_R   g1448( .A1 (n1454), .A2 (n1403), .B (n1455), .Y (y478) );
  AO21x1_ASAP7_75t_R   g1449( .A1 (n16), .A2 (n15), .B (x0), .Y (n1457) );
  INVx1_ASAP7_75t_R    g1450( .A (n1457), .Y (n1458) );
  AO32x1_ASAP7_75t_R   g1451( .A1 (n740), .A2 (n1458), .A3 (n776), .B1 (n665), .B2 (x0), .Y (y479) );
  NAND2x1_ASAP7_75t_R  g1452( .A (n15), .B (n1092), .Y (n1460) );
  AND3x1_ASAP7_75t_R   g1453( .A (n1460), .B (n1246), .C (n1247), .Y (y480) );
  INVx1_ASAP7_75t_R    g1454( .A (n67), .Y (n1462) );
  OA21x2_ASAP7_75t_R   g1455( .A1 (n1462), .A2 (n761), .B (x5), .Y (n1463) );
  AND3x1_ASAP7_75t_R   g1456( .A (n762), .B (n14), .C (y2079), .Y (n1464) );
  NOR2x1_ASAP7_75t_R   g1457( .A (n1463), .B (n1464), .Y (y481) );
  AO21x1_ASAP7_75t_R   g1458( .A1 (n15), .A2 (x5), .B (x0), .Y (n1466) );
  AO21x1_ASAP7_75t_R   g1459( .A1 (n16), .A2 (n1466), .B (n1208), .Y (n1467) );
  INVx1_ASAP7_75t_R    g1460( .A (n1467), .Y (y482) );
  INVx1_ASAP7_75t_R    g1461( .A (n276), .Y (n1469) );
  AO21x1_ASAP7_75t_R   g1462( .A1 (n15), .A2 (x3), .B (x1), .Y (n1470) );
  INVx1_ASAP7_75t_R    g1463( .A (n1470), .Y (n1471) );
  OR3x1_ASAP7_75t_R    g1464( .A (n45), .B (n16), .C (n12), .Y (n1472) );
  INVx1_ASAP7_75t_R    g1465( .A (n1472), .Y (y2220) );
  AO21x1_ASAP7_75t_R   g1466( .A1 (n1469), .A2 (n1471), .B (y2220), .Y (y483) );
  AO21x1_ASAP7_75t_R   g1467( .A1 (y9), .A2 (n45), .B (n143), .Y (n1475) );
  AO21x1_ASAP7_75t_R   g1468( .A1 (x2), .A2 (n1253), .B (n1475), .Y (y484) );
  AND3x1_ASAP7_75t_R   g1469( .A (n12), .B (x3), .C (x2), .Y (n1477) );
  AO21x1_ASAP7_75t_R   g1470( .A1 (n17), .A2 (n15), .B (n1477), .Y (n1478) );
  AO21x1_ASAP7_75t_R   g1471( .A1 (n1478), .A2 (n16), .B (n143), .Y (y485) );
  AO21x1_ASAP7_75t_R   g1472( .A1 (n16), .A2 (x3), .B (x0), .Y (n1480) );
  OA21x2_ASAP7_75t_R   g1473( .A1 (n747), .A2 (n45), .B (n1480), .Y (y486) );
  AO21x1_ASAP7_75t_R   g1474( .A1 (n17), .A2 (x2), .B (x1), .Y (n1482) );
  INVx1_ASAP7_75t_R    g1475( .A (n1482), .Y (n1483) );
  AO21x1_ASAP7_75t_R   g1476( .A1 (n15), .A2 (x3), .B (x0), .Y (n1484) );
  INVx1_ASAP7_75t_R    g1477( .A (n1484), .Y (n1485) );
  AO21x1_ASAP7_75t_R   g1478( .A1 (n1483), .A2 (n1485), .B (n143), .Y (y487) );
  OR3x1_ASAP7_75t_R    g1479( .A (n272), .B (y2079), .C (n227), .Y (y488) );
  AO21x1_ASAP7_75t_R   g1480( .A1 (x1), .A2 (x0), .B (y2079), .Y (y2813) );
  NAND2x1_ASAP7_75t_R  g1481( .A (n15), .B (y2813), .Y (n1489) );
  AO21x1_ASAP7_75t_R   g1482( .A1 (n90), .A2 (n219), .B (n15), .Y (n1490) );
  AO21x1_ASAP7_75t_R   g1483( .A1 (n1489), .A2 (n1490), .B (y2093), .Y (y489) );
  AO21x1_ASAP7_75t_R   g1484( .A1 (n12), .A2 (x5), .B (n15), .Y (n1492) );
  AO221x2_ASAP7_75t_R  g1485( .A1 (n1426), .A2 (n1492), .B1 (x2), .B2 (n989), .C (y2196), .Y (y490) );
  OR3x1_ASAP7_75t_R    g1486( .A (n225), .B (n262), .C (y2093), .Y (y491) );
  AND3x1_ASAP7_75t_R   g1487( .A (x0), .B (x2), .C (x5), .Y (n1495) );
  AND2x2_ASAP7_75t_R   g1488( .A (y25), .B (x5), .Y (n1496) );
  OAI21x1_ASAP7_75t_R  g1489( .A1 (n1496), .A2 (n854), .B (n52), .Y (n1497) );
  AO21x1_ASAP7_75t_R   g1490( .A1 (x1), .A2 (n1495), .B (n1497), .Y (y492) );
  AND3x1_ASAP7_75t_R   g1491( .A (y3293), .B (n523), .C (x0), .Y (n1499) );
  NOR2x1_ASAP7_75t_R   g1492( .A (n410), .B (n1499), .Y (y493) );
  AND3x1_ASAP7_75t_R   g1493( .A (n144), .B (n56), .C (x5), .Y (n1501) );
  AO21x1_ASAP7_75t_R   g1494( .A1 (y2079), .A2 (x0), .B (x2), .Y (n1502) );
  AND3x1_ASAP7_75t_R   g1495( .A (y3852), .B (n1502), .C (x1), .Y (n1503) );
  OR3x1_ASAP7_75t_R    g1496( .A (n1501), .B (n1503), .C (y2196), .Y (y494) );
  AO21x1_ASAP7_75t_R   g1497( .A1 (n15), .A2 (x5), .B (n227), .Y (n1505) );
  INVx1_ASAP7_75t_R    g1498( .A (y2770), .Y (n1506) );
  AND3x1_ASAP7_75t_R   g1499( .A (y2770), .B (n228), .C (n97), .Y (y3001) );
  AO21x1_ASAP7_75t_R   g1500( .A1 (n1505), .A2 (n1506), .B (y3001), .Y (y495) );
  INVx1_ASAP7_75t_R    g1501( .A (n65), .Y (n1509) );
  AO21x1_ASAP7_75t_R   g1502( .A1 (x2), .A2 (x1), .B (y2079), .Y (n1510) );
  AND3x1_ASAP7_75t_R   g1503( .A (n1469), .B (n1426), .C (x5), .Y (n1511) );
  AO21x1_ASAP7_75t_R   g1504( .A1 (n1509), .A2 (n1510), .B (n1511), .Y (y496) );
  AO21x1_ASAP7_75t_R   g1505( .A1 (n63), .A2 (n64), .B (n12), .Y (n1513) );
  NOR2x1_ASAP7_75t_R   g1506( .A (y2079), .B (n1513), .Y (n1514) );
  INVx1_ASAP7_75t_R    g1507( .A (n1514), .Y (n1515) );
  AND3x1_ASAP7_75t_R   g1508( .A (n1515), .B (n86), .C (n93), .Y (y497) );
  AND3x1_ASAP7_75t_R   g1509( .A (n244), .B (n746), .C (x1), .Y (n1517) );
  NOR2x1_ASAP7_75t_R   g1510( .A (n276), .B (n497), .Y (n1518) );
  OR3x1_ASAP7_75t_R    g1511( .A (n1517), .B (n1518), .C (y2196), .Y (y498) );
  OA33x2_ASAP7_75t_R   g1512( .A1 (n1261), .A2 (n993), .A3 (n798), .B1 (y2079), .B2 (n83), .B3 (n12), .Y (y499) );
  OR3x1_ASAP7_75t_R    g1513( .A (n13), .B (y2079), .C (n12), .Y (n1521) );
  NAND2x1_ASAP7_75t_R  g1514( .A (n12), .B (n1510), .Y (n1522) );
  AO21x1_ASAP7_75t_R   g1515( .A1 (n1521), .A2 (n1522), .B (n51), .Y (y500) );
  AO32x1_ASAP7_75t_R   g1516( .A1 (n740), .A2 (n1450), .A3 (n12), .B1 (x0), .B2 (n1336), .Y (y501) );
  INVx1_ASAP7_75t_R    g1517( .A (n1522), .Y (n1525) );
  NOR2x1_ASAP7_75t_R   g1518( .A (n1525), .B (n1514), .Y (y502) );
  INVx1_ASAP7_75t_R    g1519( .A (y25), .Y (n1527) );
  AO21x1_ASAP7_75t_R   g1520( .A1 (n15), .A2 (n16), .B (x5), .Y (n1528) );
  AO21x1_ASAP7_75t_R   g1521( .A1 (y2079), .A2 (x1), .B (x2), .Y (n1529) );
  AND2x2_ASAP7_75t_R   g1522( .A (n1529), .B (x0), .Y (n1530) );
  AO21x1_ASAP7_75t_R   g1523( .A1 (n1530), .A2 (n497), .B (n53), .Y (y2490) );
  AO21x1_ASAP7_75t_R   g1524( .A1 (n1527), .A2 (n1528), .B (y2490), .Y (y503) );
  AND2x2_ASAP7_75t_R   g1525( .A (n1336), .B (x0), .Y (y773) );
  AO21x1_ASAP7_75t_R   g1526( .A1 (n97), .A2 (y773), .B (n1501), .Y (y504) );
  NAND2x1_ASAP7_75t_R  g1527( .A (n97), .B (n64), .Y (n1535) );
  AO21x1_ASAP7_75t_R   g1528( .A1 (n16), .A2 (x2), .B (n12), .Y (n1536) );
  AND3x1_ASAP7_75t_R   g1529( .A (n15), .B (x5), .C (x1), .Y (n1537) );
  NOR2x1_ASAP7_75t_R   g1530( .A (n1536), .B (n1537), .Y (y1084) );
  AO21x1_ASAP7_75t_R   g1531( .A1 (n12), .A2 (n1535), .B (y1084), .Y (y505) );
  OR3x1_ASAP7_75t_R    g1532( .A (y863), .B (y2079), .C (x2), .Y (n1540) );
  INVx1_ASAP7_75t_R    g1533( .A (n1540), .Y (n1541) );
  AO21x1_ASAP7_75t_R   g1534( .A1 (n15), .A2 (x5), .B (n12), .Y (n1542) );
  NOR2x1_ASAP7_75t_R   g1535( .A (n16), .B (n1542), .Y (y2163) );
  OR3x1_ASAP7_75t_R    g1536( .A (n1541), .B (y2163), .C (n227), .Y (y506) );
  INVx1_ASAP7_75t_R    g1537( .A (n90), .Y (n1545) );
  AO21x1_ASAP7_75t_R   g1538( .A1 (n16), .A2 (x3), .B (x2), .Y (n1546) );
  OR3x1_ASAP7_75t_R    g1539( .A (n1545), .B (n1208), .C (n1546), .Y (n1547) );
  AND2x2_ASAP7_75t_R   g1540( .A (n1547), .B (n1490), .Y (y507) );
  AND3x1_ASAP7_75t_R   g1541( .A (n15), .B (x3), .C (x0), .Y (n1549) );
  INVx1_ASAP7_75t_R    g1542( .A (n1549), .Y (n1550) );
  AO21x1_ASAP7_75t_R   g1543( .A1 (n1550), .A2 (n244), .B (n16), .Y (n1551) );
  OA21x2_ASAP7_75t_R   g1544( .A1 (n1032), .A2 (n851), .B (n1551), .Y (y508) );
  AND3x1_ASAP7_75t_R   g1545( .A (n15), .B (x3), .C (x1), .Y (n1553) );
  INVx1_ASAP7_75t_R    g1546( .A (n1553), .Y (n1554) );
  AO21x1_ASAP7_75t_R   g1547( .A1 (n1554), .A2 (n64), .B (n12), .Y (n1555) );
  NAND2x1_ASAP7_75t_R  g1548( .A (n12), .B (n153), .Y (n1556) );
  AND2x2_ASAP7_75t_R   g1549( .A (n1555), .B (n1556), .Y (y509) );
  AND3x1_ASAP7_75t_R   g1550( .A (n12), .B (n15), .C (x3), .Y (n1558) );
  AO21x1_ASAP7_75t_R   g1551( .A1 (n72), .A2 (x0), .B (n1558), .Y (n1559) );
  AO21x1_ASAP7_75t_R   g1552( .A1 (x3), .A2 (n15), .B (n90), .Y (n1560) );
  OA21x2_ASAP7_75t_R   g1553( .A1 (n1559), .A2 (n1483), .B (n1560), .Y (y510) );
  AO21x1_ASAP7_75t_R   g1554( .A1 (n244), .A2 (n746), .B (n16), .Y (n1562) );
  OA21x2_ASAP7_75t_R   g1555( .A1 (n1032), .A2 (n851), .B (n1562), .Y (y511) );
  INVx1_ASAP7_75t_R    g1556( .A (n1536), .Y (n1564) );
  INVx1_ASAP7_75t_R    g1557( .A (n161), .Y (n1565) );
  AO21x1_ASAP7_75t_R   g1558( .A1 (n63), .A2 (n1564), .B (n1565), .Y (y512) );
  AO21x1_ASAP7_75t_R   g1559( .A1 (x3), .A2 (x2), .B (y863), .Y (n1567) );
  INVx1_ASAP7_75t_R    g1560( .A (n1567), .Y (n1568) );
  AO21x1_ASAP7_75t_R   g1561( .A1 (n16), .A2 (n12), .B (n81), .Y (n1569) );
  AND3x1_ASAP7_75t_R   g1562( .A (n103), .B (x3), .C (x0), .Y (n1570) );
  OR3x1_ASAP7_75t_R    g1563( .A (n1568), .B (n1569), .C (n1570), .Y (y513) );
  INVx1_ASAP7_75t_R    g1564( .A (n81), .Y (n1572) );
  AND3x1_ASAP7_75t_R   g1565( .A (y9), .B (n137), .C (n72), .Y (n1573) );
  AO21x1_ASAP7_75t_R   g1566( .A1 (n144), .A2 (n1572), .B (n1573), .Y (n1574) );
  NOR2x1_ASAP7_75t_R   g1567( .A (n17), .B (n1490), .Y (n1575) );
  INVx1_ASAP7_75t_R    g1568( .A (n1575), .Y (n1576) );
  NAND2x1_ASAP7_75t_R  g1569( .A (n1574), .B (n1576), .Y (n1577) );
  INVx1_ASAP7_75t_R    g1570( .A (n1577), .Y (y515) );
  AO32x1_ASAP7_75t_R   g1571( .A1 (n488), .A2 (x2), .A3 (n219), .B1 (n271), .B2 (y6), .Y (n1579) );
  AO21x1_ASAP7_75t_R   g1572( .A1 (y2079), .A2 (n228), .B (n1579), .Y (y516) );
  NOR2x1_ASAP7_75t_R   g1573( .A (y2079), .B (n1562), .Y (n1581) );
  INVx1_ASAP7_75t_R    g1574( .A (n1581), .Y (n1582) );
  INVx1_ASAP7_75t_R    g1575( .A (n1495), .Y (n1583) );
  AO21x1_ASAP7_75t_R   g1576( .A1 (n1583), .A2 (n751), .B (x1), .Y (n1584) );
  AND2x2_ASAP7_75t_R   g1577( .A (n1582), .B (n1584), .Y (y517) );
  AO21x1_ASAP7_75t_R   g1578( .A1 (n63), .A2 (n64), .B (y2079), .Y (n1586) );
  NOR2x1_ASAP7_75t_R   g1579( .A (x0), .B (n1586), .Y (n1587) );
  AO21x1_ASAP7_75t_R   g1580( .A1 (n63), .A2 (n64), .B (x0), .Y (y1116) );
  AND2x2_ASAP7_75t_R   g1581( .A (y1116), .B (y2079), .Y (y2787) );
  AO21x1_ASAP7_75t_R   g1582( .A1 (x1), .A2 (n15), .B (n1536), .Y (n1590) );
  INVx1_ASAP7_75t_R    g1583( .A (n1590), .Y (y2259) );
  OR3x1_ASAP7_75t_R    g1584( .A (n1587), .B (y2787), .C (y2259), .Y (y518) );
  OA21x2_ASAP7_75t_R   g1585( .A1 (x0), .A2 (n801), .B (n737), .Y (y519) );
  AO21x1_ASAP7_75t_R   g1586( .A1 (n90), .A2 (n219), .B (x2), .Y (n1594) );
  NAND2x1_ASAP7_75t_R  g1587( .A (x5), .B (n1594), .Y (n1595) );
  AND3x1_ASAP7_75t_R   g1588( .A (n90), .B (n219), .C (x2), .Y (n1596) );
  AND2x2_ASAP7_75t_R   g1589( .A (n174), .B (n1312), .Y (n1597) );
  INVx1_ASAP7_75t_R    g1590( .A (n1597), .Y (n1598) );
  OA21x2_ASAP7_75t_R   g1591( .A1 (n1595), .A2 (n1596), .B (n1598), .Y (y520) );
  AO21x1_ASAP7_75t_R   g1592( .A1 (n12), .A2 (x2), .B (x5), .Y (n1600) );
  INVx1_ASAP7_75t_R    g1593( .A (n1600), .Y (n1601) );
  AO21x1_ASAP7_75t_R   g1594( .A1 (n1509), .A2 (n1513), .B (n1601), .Y (y521) );
  AO21x1_ASAP7_75t_R   g1595( .A1 (n16), .A2 (x0), .B (x5), .Y (n1603) );
  INVx1_ASAP7_75t_R    g1596( .A (n1603), .Y (n1604) );
  OR4x2_ASAP7_75t_R    g1597( .A (n1208), .B (n1604), .C (n1245), .D (x2), .Y (n1605) );
  AO21x1_ASAP7_75t_R   g1598( .A1 (n1246), .A2 (n219), .B (n15), .Y (n1606) );
  AND2x2_ASAP7_75t_R   g1599( .A (n1605), .B (n1606), .Y (y522) );
  INVx1_ASAP7_75t_R    g1600( .A (n1380), .Y (n1608) );
  AO21x1_ASAP7_75t_R   g1601( .A1 (n15), .A2 (n1608), .B (n1596), .Y (y523) );
  AO21x1_ASAP7_75t_R   g1602( .A1 (n12), .A2 (n497), .B (n1245), .Y (n1610) );
  INVx1_ASAP7_75t_R    g1603( .A (n1610), .Y (y1553) );
  OA22x2_ASAP7_75t_R   g1604( .A1 (n15), .A2 (y1553), .B1 (n97), .B2 (n1610), .Y (y524) );
  INVx1_ASAP7_75t_R    g1605( .A (n113), .Y (n1613) );
  AO21x1_ASAP7_75t_R   g1606( .A1 (n64), .A2 (n63), .B (y2079), .Y (n1614) );
  AND2x2_ASAP7_75t_R   g1607( .A (n1614), .B (x0), .Y (n1615) );
  AO21x1_ASAP7_75t_R   g1608( .A1 (n753), .A2 (n1613), .B (n1615), .Y (y525) );
  AND2x2_ASAP7_75t_R   g1609( .A (n455), .B (n84), .Y (n1617) );
  AO21x1_ASAP7_75t_R   g1610( .A1 (x4), .A2 (x5), .B (n145), .Y (n1618) );
  INVx1_ASAP7_75t_R    g1611( .A (n1618), .Y (n1619) );
  AO21x1_ASAP7_75t_R   g1612( .A1 (n388), .A2 (n28), .B (x3), .Y (n1620) );
  OA21x2_ASAP7_75t_R   g1613( .A1 (n1617), .A2 (n1619), .B (n1620), .Y (y526) );
  NOR2x1_ASAP7_75t_R   g1614( .A (n606), .B (n410), .Y (y527) );
  AND3x1_ASAP7_75t_R   g1615( .A (n16), .B (x2), .C (x5), .Y (n1623) );
  INVx1_ASAP7_75t_R    g1616( .A (n1623), .Y (n1624) );
  AO21x1_ASAP7_75t_R   g1617( .A1 (n15), .A2 (n497), .B (n1623), .Y (n1625) );
  AO32x1_ASAP7_75t_R   g1618( .A1 (n1624), .A2 (n750), .A3 (x0), .B1 (n1092), .B2 (n1625), .Y (y528) );
  AO21x1_ASAP7_75t_R   g1619( .A1 (n1510), .A2 (x0), .B (n51), .Y (n1627) );
  AO21x1_ASAP7_75t_R   g1620( .A1 (y19), .A2 (n1627), .B (n1587), .Y (y529) );
  INVx1_ASAP7_75t_R    g1621( .A (n1586), .Y (n1629) );
  AND2x2_ASAP7_75t_R   g1622( .A (n1586), .B (x0), .Y (y1067) );
  AO21x1_ASAP7_75t_R   g1623( .A1 (n12), .A2 (n1629), .B (y1067), .Y (y530) );
  AND3x1_ASAP7_75t_R   g1624( .A (n178), .B (n1528), .C (n14), .Y (n1632) );
  NOR2x1_ASAP7_75t_R   g1625( .A (n12), .B (n1632), .Y (y1069) );
  AO21x1_ASAP7_75t_R   g1626( .A1 (n12), .A2 (n1632), .B (y1069), .Y (y531) );
  AO21x1_ASAP7_75t_R   g1627( .A1 (n12), .A2 (n16), .B (x2), .Y (n1635) );
  INVx1_ASAP7_75t_R    g1628( .A (n1635), .Y (n1636) );
  AND3x1_ASAP7_75t_R   g1629( .A (n97), .B (n219), .C (n90), .Y (n1637) );
  AO21x1_ASAP7_75t_R   g1630( .A1 (n988), .A2 (n1636), .B (n1637), .Y (y532) );
  AO21x1_ASAP7_75t_R   g1631( .A1 (n544), .A2 (n15), .B (x0), .Y (n1639) );
  INVx1_ASAP7_75t_R    g1632( .A (n1537), .Y (n1640) );
  AO21x1_ASAP7_75t_R   g1633( .A1 (n1640), .A2 (n64), .B (n12), .Y (n1641) );
  OA21x2_ASAP7_75t_R   g1634( .A1 (n1262), .A2 (n1639), .B (n1641), .Y (y533) );
  INVx1_ASAP7_75t_R    g1635( .A (n99), .Y (n1643) );
  AND3x1_ASAP7_75t_R   g1636( .A (n16), .B (n15), .C (x5), .Y (n1644) );
  OR3x1_ASAP7_75t_R    g1637( .A (n798), .B (n1643), .C (n1644), .Y (y534) );
  INVx1_ASAP7_75t_R    g1638( .A (n97), .Y (n1646) );
  AND3x1_ASAP7_75t_R   g1639( .A (n97), .B (n90), .C (n219), .Y (n1647) );
  AO21x1_ASAP7_75t_R   g1640( .A1 (n221), .A2 (n1646), .B (n1647), .Y (y535) );
  AND3x1_ASAP7_75t_R   g1641( .A (n241), .B (n16), .C (x5), .Y (n1649) );
  AO21x1_ASAP7_75t_R   g1642( .A1 (n1540), .A2 (n228), .B (n1649), .Y (y536) );
  NAND2x1_ASAP7_75t_R  g1643( .A (n15), .B (n1242), .Y (n1651) );
  XOR2x2_ASAP7_75t_R   g1644( .A (n221), .B (n1651), .Y (y537) );
  INVx1_ASAP7_75t_R    g1645( .A (n1490), .Y (n1653) );
  NOR2x1_ASAP7_75t_R   g1646( .A (n1234), .B (n1653), .Y (y538) );
  AO32x1_ASAP7_75t_R   g1647( .A1 (n12), .A2 (y3293), .A3 (x1), .B1 (y1894), .B2 (n469), .Y (y539) );
  AO21x1_ASAP7_75t_R   g1648( .A1 (n12), .A2 (x3), .B (x1), .Y (n1656) );
  INVx1_ASAP7_75t_R    g1649( .A (n184), .Y (n1657) );
  AO32x1_ASAP7_75t_R   g1650( .A1 (n72), .A2 (n219), .A3 (n1656), .B1 (n271), .B2 (n1657), .Y (y540) );
  AO21x1_ASAP7_75t_R   g1651( .A1 (n64), .A2 (n63), .B (n17), .Y (n1659) );
  INVx1_ASAP7_75t_R    g1652( .A (n1659), .Y (n1660) );
  NOR2x1_ASAP7_75t_R   g1653( .A (n1536), .B (n1553), .Y (n1661) );
  AO21x1_ASAP7_75t_R   g1654( .A1 (n12), .A2 (n1660), .B (n1661), .Y (y541) );
  AO21x1_ASAP7_75t_R   g1655( .A1 (n241), .A2 (n993), .B (y58), .Y (y542) );
  AO21x1_ASAP7_75t_R   g1656( .A1 (n244), .A2 (n746), .B (n17), .Y (n1664) );
  NOR2x1_ASAP7_75t_R   g1657( .A (x1), .B (n1664), .Y (n1665) );
  AO21x1_ASAP7_75t_R   g1658( .A1 (n1559), .A2 (x1), .B (n1665), .Y (y543) );
  NAND2x1_ASAP7_75t_R  g1659( .A (n1656), .B (n219), .Y (n1667) );
  INVx1_ASAP7_75t_R    g1660( .A (n1667), .Y (n1668) );
  INVx1_ASAP7_75t_R    g1661( .A (n1594), .Y (n1669) );
  AO21x1_ASAP7_75t_R   g1662( .A1 (x2), .A2 (n1668), .B (n1669), .Y (y544) );
  AO21x1_ASAP7_75t_R   g1663( .A1 (n63), .A2 (n64), .B (n17), .Y (n1671) );
  INVx1_ASAP7_75t_R    g1664( .A (n1671), .Y (n1672) );
  AO21x1_ASAP7_75t_R   g1665( .A1 (n1672), .A2 (n12), .B (y2259), .Y (y545) );
  NAND2x1_ASAP7_75t_R  g1666( .A (x0), .B (n763), .Y (n1674) );
  INVx1_ASAP7_75t_R    g1667( .A (n1674), .Y (n1675) );
  INVx1_ASAP7_75t_R    g1668( .A (n694), .Y (n1676) );
  AO32x1_ASAP7_75t_R   g1669( .A1 (n63), .A2 (n64), .A3 (n1675), .B1 (n1676), .B2 (n1674), .Y (y546) );
  INVx1_ASAP7_75t_R    g1670( .A (n1480), .Y (n1678) );
  NOR2x1_ASAP7_75t_R   g1671( .A (x3), .B (n43), .Y (n1679) );
  NOR2x1_ASAP7_75t_R   g1672( .A (x2), .B (n1679), .Y (n1680) );
  OA33x2_ASAP7_75t_R   g1673( .A1 (x2), .A2 (n1678), .A3 (n1545), .B1 (n1253), .B2 (n1680), .B3 (n143), .Y (y547) );
  AND3x1_ASAP7_75t_R   g1674( .A (x1), .B (x0), .C (x3), .Y (n1682) );
  INVx1_ASAP7_75t_R    g1675( .A (n1682), .Y (n1683) );
  AO21x1_ASAP7_75t_R   g1676( .A1 (n1683), .A2 (n228), .B (n15), .Y (n1684) );
  OR3x1_ASAP7_75t_R    g1677( .A (n1682), .B (n227), .C (x2), .Y (n1685) );
  AND3x1_ASAP7_75t_R   g1678( .A (n1684), .B (n1685), .C (n260), .Y (n1686) );
  INVx1_ASAP7_75t_R    g1679( .A (n1686), .Y (y548) );
  AO21x1_ASAP7_75t_R   g1680( .A1 (x0), .A2 (n243), .B (n227), .Y (n1688) );
  NAND2x1_ASAP7_75t_R  g1681( .A (x2), .B (n260), .Y (n1689) );
  AO21x1_ASAP7_75t_R   g1682( .A1 (n1683), .A2 (n228), .B (x2), .Y (n1690) );
  OA21x2_ASAP7_75t_R   g1683( .A1 (n1688), .A2 (n1689), .B (n1690), .Y (y549) );
  AND3x1_ASAP7_75t_R   g1684( .A (n90), .B (n219), .C (x3), .Y (n1692) );
  INVx1_ASAP7_75t_R    g1685( .A (n1596), .Y (n1693) );
  AO21x1_ASAP7_75t_R   g1686( .A1 (n1693), .A2 (n17), .B (n1669), .Y (n1694) );
  AO21x1_ASAP7_75t_R   g1687( .A1 (x2), .A2 (n1692), .B (n1694), .Y (y550) );
  AND3x1_ASAP7_75t_R   g1688( .A (n17), .B (n15), .C (x1), .Y (n1696) );
  INVx1_ASAP7_75t_R    g1689( .A (n1696), .Y (n1697) );
  AO21x1_ASAP7_75t_R   g1690( .A1 (x3), .A2 (x2), .B (n12), .Y (n1698) );
  INVx1_ASAP7_75t_R    g1691( .A (n1477), .Y (n1699) );
  AO21x1_ASAP7_75t_R   g1692( .A1 (n77), .A2 (x0), .B (n1477), .Y (n1700) );
  AO32x1_ASAP7_75t_R   g1693( .A1 (n1698), .A2 (n1699), .A3 (n16), .B1 (x1), .B2 (n1700), .Y (n1701) );
  NAND2x1_ASAP7_75t_R  g1694( .A (n1697), .B (n1701), .Y (y551) );
  OR3x1_ASAP7_75t_R    g1695( .A (n128), .B (n12), .C (x3), .Y (n1703) );
  AND2x2_ASAP7_75t_R   g1696( .A (n1703), .B (n84), .Y (n1704) );
  INVx1_ASAP7_75t_R    g1697( .A (n1703), .Y (n1705) );
  OA33x2_ASAP7_75t_R   g1698( .A1 (n1261), .A2 (n1262), .A3 (n1704), .B1 (n1705), .B2 (n694), .B3 (n1032), .Y (y552) );
  AO21x1_ASAP7_75t_R   g1699( .A1 (n16), .A2 (n12), .B (x4), .Y (n1707) );
  INVx1_ASAP7_75t_R    g1700( .A (n1707), .Y (n1708) );
  OR3x1_ASAP7_75t_R    g1701( .A (y3758), .B (n1708), .C (y863), .Y (y553) );
  AO21x1_ASAP7_75t_R   g1702( .A1 (n469), .A2 (y3293), .B (n143), .Y (y554) );
  OR3x1_ASAP7_75t_R    g1703( .A (n529), .B (n29), .C (n977), .Y (y556) );
  AO21x1_ASAP7_75t_R   g1704( .A1 (n244), .A2 (n746), .B (x5), .Y (n1712) );
  AND3x1_ASAP7_75t_R   g1705( .A (n1712), .B (n1440), .C (n219), .Y (y557) );
  OR3x1_ASAP7_75t_R    g1706( .A (n529), .B (n29), .C (y863), .Y (y558) );
  AO21x1_ASAP7_75t_R   g1707( .A1 (n64), .A2 (y2079), .B (n58), .Y (n1715) );
  AND2x2_ASAP7_75t_R   g1708( .A (n1715), .B (n784), .Y (y559) );
  INVx1_ASAP7_75t_R    g1709( .A (y3428), .Y (n1717) );
  OR3x1_ASAP7_75t_R    g1710( .A (y863), .B (n22), .C (y2079), .Y (n1718) );
  AND2x2_ASAP7_75t_R   g1711( .A (n1717), .B (n1718), .Y (y560) );
  OR3x1_ASAP7_75t_R    g1712( .A (n143), .B (n22), .C (y2079), .Y (n1720) );
  AND2x2_ASAP7_75t_R   g1713( .A (n469), .B (n1720), .Y (y561) );
  AO21x1_ASAP7_75t_R   g1714( .A1 (y2813), .A2 (x4), .B (n29), .Y (y562) );
  AO21x1_ASAP7_75t_R   g1715( .A1 (n299), .A2 (x1), .B (y1281), .Y (y563) );
  NAND2x1_ASAP7_75t_R  g1716( .A (n388), .B (n310), .Y (y1300) );
  AO21x1_ASAP7_75t_R   g1717( .A1 (n544), .A2 (n299), .B (y1300), .Y (y564) );
  OR3x1_ASAP7_75t_R    g1718( .A (n43), .B (y2079), .C (x4), .Y (n1726) );
  INVx1_ASAP7_75t_R    g1719( .A (n1726), .Y (n1727) );
  OR3x1_ASAP7_75t_R    g1720( .A (n1727), .B (n143), .C (n529), .Y (y565) );
  AO21x1_ASAP7_75t_R   g1721( .A1 (x1), .A2 (x0), .B (x4), .Y (n1729) );
  INVx1_ASAP7_75t_R    g1722( .A (n1729), .Y (n1730) );
  AO21x1_ASAP7_75t_R   g1723( .A1 (x0), .A2 (n544), .B (n1730), .Y (n1731) );
  AO21x1_ASAP7_75t_R   g1724( .A1 (n1731), .A2 (n228), .B (n529), .Y (y566) );
  AO21x1_ASAP7_75t_R   g1725( .A1 (y3852), .A2 (n125), .B (n1278), .Y (y567) );
  OA21x2_ASAP7_75t_R   g1726( .A1 (n1454), .A2 (n1403), .B (y3852), .Y (y568) );
  AND2x2_ASAP7_75t_R   g1727( .A (y563), .B (n453), .Y (y569) );
  AO21x1_ASAP7_75t_R   g1728( .A1 (y9), .A2 (y3293), .B (n143), .Y (y570) );
  AND3x1_ASAP7_75t_R   g1729( .A (n1240), .B (n1707), .C (y2079), .Y (n1737) );
  OR3x1_ASAP7_75t_R    g1730( .A (n227), .B (y2079), .C (x4), .Y (n1738) );
  INVx1_ASAP7_75t_R    g1731( .A (n1738), .Y (n1739) );
  OR3x1_ASAP7_75t_R    g1732( .A (n1737), .B (n1739), .C (y863), .Y (y571) );
  AND2x2_ASAP7_75t_R   g1733( .A (y558), .B (n228), .Y (y572) );
  OR3x1_ASAP7_75t_R    g1734( .A (y2466), .B (x0), .C (x1), .Y (n1742) );
  INVx1_ASAP7_75t_R    g1735( .A (n34), .Y (n1743) );
  OR3x1_ASAP7_75t_R    g1736( .A (y2466), .B (n12), .C (n16), .Y (n1744) );
  INVx1_ASAP7_75t_R    g1737( .A (n1744), .Y (n1745) );
  AO21x1_ASAP7_75t_R   g1738( .A1 (n1742), .A2 (n1743), .B (n1745), .Y (y573) );
  AO21x1_ASAP7_75t_R   g1739( .A1 (n12), .A2 (x4), .B (n16), .Y (n1747) );
  INVx1_ASAP7_75t_R    g1740( .A (n1747), .Y (n1748) );
  AO21x1_ASAP7_75t_R   g1741( .A1 (n22), .A2 (y3852), .B (n1748), .Y (n1749) );
  OR3x1_ASAP7_75t_R    g1742( .A (n43), .B (n22), .C (x5), .Y (n1750) );
  INVx1_ASAP7_75t_R    g1743( .A (n1750), .Y (n1751) );
  AO21x1_ASAP7_75t_R   g1744( .A1 (n1749), .A2 (n1106), .B (n1751), .Y (y574) );
  AO21x1_ASAP7_75t_R   g1745( .A1 (y2079), .A2 (n108), .B (y1081), .Y (y575) );
  AND2x2_ASAP7_75t_R   g1746( .A (y562), .B (n228), .Y (y576) );
  AO21x1_ASAP7_75t_R   g1747( .A1 (n28), .A2 (n352), .B (x1), .Y (n1755) );
  AND2x2_ASAP7_75t_R   g1748( .A (n1755), .B (y104), .Y (y577) );
  AND3x1_ASAP7_75t_R   g1749( .A (n363), .B (n22), .C (n16), .Y (n1757) );
  INVx1_ASAP7_75t_R    g1750( .A (n1757), .Y (n1758) );
  OR3x1_ASAP7_75t_R    g1751( .A (n527), .B (y2079), .C (n143), .Y (y2432) );
  AND2x2_ASAP7_75t_R   g1752( .A (n1758), .B (y2432), .Y (y578) );
  AND2x2_ASAP7_75t_R   g1753( .A (n445), .B (y2432), .Y (y579) );
  AO21x1_ASAP7_75t_R   g1754( .A1 (y2079), .A2 (x4), .B (n527), .Y (n1762) );
  AO21x1_ASAP7_75t_R   g1755( .A1 (x0), .A2 (x1), .B (n1762), .Y (y580) );
  OA21x2_ASAP7_75t_R   g1756( .A1 (n993), .A2 (n604), .B (n1191), .Y (y581) );
  NAND2x1_ASAP7_75t_R  g1757( .A (n824), .B (n797), .Y (y582) );
  NAND2x1_ASAP7_75t_R  g1758( .A (n17), .B (n174), .Y (n1766) );
  NAND2x1_ASAP7_75t_R  g1759( .A (n747), .B (n219), .Y (n1767) );
  INVx1_ASAP7_75t_R    g1760( .A (n1767), .Y (n1768) );
  XNOR2x2_ASAP7_75t_R  g1761( .A (n1766), .B (n1768), .Y (y583) );
  NOR2x1_ASAP7_75t_R   g1762( .A (x1), .B (n473), .Y (n1770) );
  OR3x1_ASAP7_75t_R    g1763( .A (n1016), .B (n1770), .C (n529), .Y (y584) );
  INVx1_ASAP7_75t_R    g1764( .A (n1644), .Y (n1772) );
  AO21x1_ASAP7_75t_R   g1765( .A1 (n1772), .A2 (x0), .B (n495), .Y (y585) );
  AND2x2_ASAP7_75t_R   g1766( .A (n466), .B (n219), .Y (n1774) );
  INVx1_ASAP7_75t_R    g1767( .A (n614), .Y (n1775) );
  AO21x1_ASAP7_75t_R   g1768( .A1 (n1774), .A2 (x5), .B (n1775), .Y (y586) );
  AO21x1_ASAP7_75t_R   g1769( .A1 (n1774), .A2 (x5), .B (n972), .Y (y587) );
  AND3x1_ASAP7_75t_R   g1770( .A (x0), .B (x1), .C (x5), .Y (n1778) );
  AO21x1_ASAP7_75t_R   g1771( .A1 (y2079), .A2 (x4), .B (n1778), .Y (n1779) );
  AO21x1_ASAP7_75t_R   g1772( .A1 (n474), .A2 (n16), .B (n1779), .Y (y588) );
  AND2x2_ASAP7_75t_R   g1773( .A (n1114), .B (n1026), .Y (y589) );
  AO21x1_ASAP7_75t_R   g1774( .A1 (x0), .A2 (x1), .B (y2079), .Y (n1782) );
  AND2x2_ASAP7_75t_R   g1775( .A (y9), .B (n1782), .Y (y741) );
  OA21x2_ASAP7_75t_R   g1776( .A1 (n527), .A2 (y741), .B (n445), .Y (y590) );
  AND2x2_ASAP7_75t_R   g1777( .A (n64), .B (n219), .Y (n1785) );
  AO21x1_ASAP7_75t_R   g1778( .A1 (x0), .A2 (n16), .B (n72), .Y (n1786) );
  NOR2x1_ASAP7_75t_R   g1779( .A (x0), .B (n1659), .Y (n1787) );
  AO21x1_ASAP7_75t_R   g1780( .A1 (n1785), .A2 (n1786), .B (n1787), .Y (y591) );
  OR3x1_ASAP7_75t_R    g1781( .A (n989), .B (n990), .C (n478), .Y (y592) );
  AO22x1_ASAP7_75t_R   g1782( .A1 (n16), .A2 (n718), .B1 (x1), .B2 (n604), .Y (y593) );
  OR3x1_ASAP7_75t_R    g1783( .A (x5), .B (x4), .C (x3), .Y (n1791) );
  AND2x2_ASAP7_75t_R   g1784( .A (y193), .B (n1791), .Y (y594) );
  AND3x1_ASAP7_75t_R   g1785( .A (n455), .B (n776), .C (n466), .Y (n1793) );
  AO21x1_ASAP7_75t_R   g1786( .A1 (n497), .A2 (x0), .B (n1793), .Y (y595) );
  AO21x1_ASAP7_75t_R   g1787( .A1 (n770), .A2 (x0), .B (n701), .Y (y596) );
  AO21x1_ASAP7_75t_R   g1788( .A1 (n529), .A2 (y9), .B (n143), .Y (n1796) );
  AO21x1_ASAP7_75t_R   g1789( .A1 (n527), .A2 (n352), .B (n1796), .Y (y597) );
  AO21x1_ASAP7_75t_R   g1790( .A1 (n352), .A2 (x1), .B (n990), .Y (n1798) );
  AO21x1_ASAP7_75t_R   g1791( .A1 (n1798), .A2 (y3852), .B (n527), .Y (y598) );
  AO21x1_ASAP7_75t_R   g1792( .A1 (n139), .A2 (n16), .B (n143), .Y (n1800) );
  AO21x1_ASAP7_75t_R   g1793( .A1 (n211), .A2 (y9), .B (n1800), .Y (y599) );
  AO21x1_ASAP7_75t_R   g1794( .A1 (n583), .A2 (n439), .B (n16), .Y (n1802) );
  NAND2x1_ASAP7_75t_R  g1795( .A (n1755), .B (n1802), .Y (y600) );
  AO32x1_ASAP7_75t_R   g1796( .A1 (n466), .A2 (n352), .A3 (n1026), .B1 (x0), .B2 (n529), .Y (y601) );
  AND3x1_ASAP7_75t_R   g1797( .A (y9), .B (n310), .C (y2079), .Y (n1805) );
  AO21x1_ASAP7_75t_R   g1798( .A1 (n1774), .A2 (x5), .B (n1805), .Y (y602) );
  AO21x1_ASAP7_75t_R   g1799( .A1 (n90), .A2 (n219), .B (y3758), .Y (y603) );
  OA21x2_ASAP7_75t_R   g1800( .A1 (x0), .A2 (n998), .B (n963), .Y (y604) );
  AO21x1_ASAP7_75t_R   g1801( .A1 (y2079), .A2 (x4), .B (y863), .Y (n1809) );
  AO21x1_ASAP7_75t_R   g1802( .A1 (x5), .A2 (n948), .B (n1809), .Y (y605) );
  AO21x1_ASAP7_75t_R   g1803( .A1 (n1774), .A2 (n352), .B (n1004), .Y (y606) );
  AND3x1_ASAP7_75t_R   g1804( .A (n1114), .B (n1026), .C (n455), .Y (y607) );
  AO21x1_ASAP7_75t_R   g1805( .A1 (y3852), .A2 (n90), .B (n527), .Y (y608) );
  AO32x1_ASAP7_75t_R   g1806( .A1 (n466), .A2 (n219), .A3 (n583), .B1 (n363), .B2 (n534), .Y (y609) );
  NAND2x1_ASAP7_75t_R  g1807( .A (n488), .B (n219), .Y (n1815) );
  OA21x2_ASAP7_75t_R   g1808( .A1 (n1815), .A2 (x2), .B (n1490), .Y (y610) );
  AND3x1_ASAP7_75t_R   g1809( .A (n12), .B (y2079), .C (x4), .Y (n1817) );
  OR3x1_ASAP7_75t_R    g1810( .A (n478), .B (n1817), .C (n143), .Y (y611) );
  AND2x2_ASAP7_75t_R   g1811( .A (y3852), .B (n90), .Y (n1819) );
  AO21x1_ASAP7_75t_R   g1812( .A1 (n1819), .A2 (n455), .B (n527), .Y (y612) );
  AND2x2_ASAP7_75t_R   g1813( .A (n1064), .B (y608), .Y (y613) );
  AND2x2_ASAP7_75t_R   g1814( .A (y608), .B (n455), .Y (y614) );
  AO21x1_ASAP7_75t_R   g1815( .A1 (x0), .A2 (x1), .B (n606), .Y (y615) );
  NOR2x1_ASAP7_75t_R   g1816( .A (n186), .B (n1541), .Y (y616) );
  AO21x1_ASAP7_75t_R   g1817( .A1 (n28), .A2 (n614), .B (x1), .Y (n1825) );
  NAND2x1_ASAP7_75t_R  g1818( .A (n144), .B (n1825), .Y (y617) );
  AND2x2_ASAP7_75t_R   g1819( .A (y3852), .B (n763), .Y (y618) );
  NOR2x1_ASAP7_75t_R   g1820( .A (n1208), .B (n1045), .Y (y619) );
  AND2x2_ASAP7_75t_R   g1821( .A (y3293), .B (n523), .Y (n1829) );
  NOR2x1_ASAP7_75t_R   g1822( .A (n436), .B (n352), .Y (n1830) );
  INVx1_ASAP7_75t_R    g1823( .A (n1830), .Y (n1831) );
  OA21x2_ASAP7_75t_R   g1824( .A1 (n143), .A2 (n1829), .B (n1831), .Y (y620) );
  AND3x1_ASAP7_75t_R   g1825( .A (n1064), .B (n1191), .C (n219), .Y (y622) );
  NAND2x1_ASAP7_75t_R  g1826( .A (x5), .B (n976), .Y (y623) );
  NAND2x1_ASAP7_75t_R  g1827( .A (n976), .B (n697), .Y (y624) );
  AO21x1_ASAP7_75t_R   g1828( .A1 (y2079), .A2 (n976), .B (n1083), .Y (y625) );
  AO21x1_ASAP7_75t_R   g1829( .A1 (y2079), .A2 (n436), .B (n977), .Y (y626) );
  INVx1_ASAP7_75t_R    g1830( .A (n211), .Y (n1838) );
  AO21x1_ASAP7_75t_R   g1831( .A1 (n15), .A2 (n17), .B (n16), .Y (n1839) );
  AO21x1_ASAP7_75t_R   g1832( .A1 (n1838), .A2 (n1839), .B (n12), .Y (n1840) );
  AO21x1_ASAP7_75t_R   g1833( .A1 (x0), .A2 (x1), .B (x3), .Y (n1841) );
  INVx1_ASAP7_75t_R    g1834( .A (n1841), .Y (n1842) );
  AND2x2_ASAP7_75t_R   g1835( .A (n56), .B (n1842), .Y (n1843) );
  INVx1_ASAP7_75t_R    g1836( .A (n1843), .Y (n1844) );
  NAND2x1_ASAP7_75t_R  g1837( .A (n1840), .B (n1844), .Y (y627) );
  AO21x1_ASAP7_75t_R   g1838( .A1 (n12), .A2 (n16), .B (x4), .Y (n1846) );
  AO21x1_ASAP7_75t_R   g1839( .A1 (y2079), .A2 (n1846), .B (n1083), .Y (y628) );
  AO21x1_ASAP7_75t_R   g1840( .A1 (n1093), .A2 (n466), .B (n1775), .Y (y629) );
  AO21x1_ASAP7_75t_R   g1841( .A1 (n1093), .A2 (n466), .B (n529), .Y (y631) );
  AND2x2_ASAP7_75t_R   g1842( .A (y623), .B (n453), .Y (y632) );
  INVx1_ASAP7_75t_R    g1843( .A (n315), .Y (n1851) );
  AO221x2_ASAP7_75t_R  g1844( .A1 (x0), .A2 (x5), .B1 (n1851), .B2 (n628), .C (n630), .Y (y634) );
  INVx1_ASAP7_75t_R    g1845( .A (n974), .Y (n1853) );
  AO21x1_ASAP7_75t_R   g1846( .A1 (n1853), .A2 (y2079), .B (n977), .Y (y635) );
  AO21x1_ASAP7_75t_R   g1847( .A1 (y2079), .A2 (n511), .B (n1184), .Y (y636) );
  AND2x2_ASAP7_75t_R   g1848( .A (n1356), .B (n228), .Y (y637) );
  AND2x2_ASAP7_75t_R   g1849( .A (n443), .B (n1114), .Y (y638) );
  AO21x1_ASAP7_75t_R   g1850( .A1 (n495), .A2 (x4), .B (x0), .Y (n1858) );
  AND2x2_ASAP7_75t_R   g1851( .A (n1858), .B (n1191), .Y (y639) );
  AND2x2_ASAP7_75t_R   g1852( .A (n1846), .B (y2079), .Y (n1860) );
  OA21x2_ASAP7_75t_R   g1853( .A1 (n1860), .A2 (n530), .B (n1114), .Y (y640) );
  NOR2x1_ASAP7_75t_R   g1854( .A (n312), .B (n310), .Y (n1862) );
  INVx1_ASAP7_75t_R    g1855( .A (n1862), .Y (n1863) );
  AND3x1_ASAP7_75t_R   g1856( .A (n1863), .B (n1114), .C (y3852), .Y (y641) );
  AO21x1_ASAP7_75t_R   g1857( .A1 (n1774), .A2 (n352), .B (n529), .Y (y642) );
  AND3x1_ASAP7_75t_R   g1858( .A (n1114), .B (n546), .C (y3852), .Y (y643) );
  AO21x1_ASAP7_75t_R   g1859( .A1 (n1774), .A2 (x5), .B (n529), .Y (y644) );
  AND2x2_ASAP7_75t_R   g1860( .A (n963), .B (y195), .Y (y645) );
  AND2x2_ASAP7_75t_R   g1861( .A (n1008), .B (y623), .Y (y646) );
  AO21x1_ASAP7_75t_R   g1862( .A1 (x2), .A2 (y2079), .B (n90), .Y (n1870) );
  AND2x2_ASAP7_75t_R   g1863( .A (n1870), .B (n219), .Y (y647) );
  AO21x1_ASAP7_75t_R   g1864( .A1 (n466), .A2 (x0), .B (n363), .Y (y648) );
  OR3x1_ASAP7_75t_R    g1865( .A (x1), .B (x3), .C (x2), .Y (n1873) );
  INVx1_ASAP7_75t_R    g1866( .A (n1873), .Y (n1874) );
  AO21x1_ASAP7_75t_R   g1867( .A1 (n883), .A2 (x0), .B (n1874), .Y (y649) );
  AND2x2_ASAP7_75t_R   g1868( .A (n1125), .B (y3852), .Y (y650) );
  AO21x1_ASAP7_75t_R   g1869( .A1 (n436), .A2 (n363), .B (n977), .Y (y651) );
  INVx1_ASAP7_75t_R    g1870( .A (n1050), .Y (n1878) );
  AO21x1_ASAP7_75t_R   g1871( .A1 (n16), .A2 (n22), .B (n12), .Y (n1879) );
  OA21x2_ASAP7_75t_R   g1872( .A1 (n1878), .A2 (n1879), .B (y3852), .Y (y652) );
  NAND2x1_ASAP7_75t_R  g1873( .A (n12), .B (n697), .Y (n1881) );
  OA21x2_ASAP7_75t_R   g1874( .A1 (n1878), .A2 (n1879), .B (n1881), .Y (y653) );
  OR3x1_ASAP7_75t_R    g1875( .A (n529), .B (n29), .C (n427), .Y (y654) );
  AO21x1_ASAP7_75t_R   g1876( .A1 (n1000), .A2 (x0), .B (n363), .Y (y655) );
  INVx1_ASAP7_75t_R    g1877( .A (n252), .Y (n1885) );
  AO21x1_ASAP7_75t_R   g1878( .A1 (x1), .A2 (x3), .B (x0), .Y (n1886) );
  INVx1_ASAP7_75t_R    g1879( .A (n1886), .Y (n1887) );
  AO221x2_ASAP7_75t_R  g1880( .A1 (n1885), .A2 (n1887), .B1 (n252), .B2 (n1886), .C (n143), .Y (y656) );
  AO21x1_ASAP7_75t_R   g1881( .A1 (n15), .A2 (x0), .B (y2079), .Y (n1889) );
  AOI22x1_ASAP7_75t_R  g1882( .A1 (n16), .A2 (n1889), .B1 (n1458), .B2 (n740), .Y (y657) );
  NAND2x1_ASAP7_75t_R  g1883( .A (y2466), .B (n219), .Y (n1891) );
  AND2x2_ASAP7_75t_R   g1884( .A (n1891), .B (y648), .Y (y658) );
  AND3x1_ASAP7_75t_R   g1885( .A (n546), .B (n968), .C (y3852), .Y (y659) );
  OR3x1_ASAP7_75t_R    g1886( .A (x2), .B (x3), .C (x1), .Y (n1894) );
  AO21x1_ASAP7_75t_R   g1887( .A1 (n13), .A2 (x3), .B (x0), .Y (y1110) );
  AND3x1_ASAP7_75t_R   g1888( .A (n43), .B (n17), .C (n15), .Y (n1896) );
  AO21x1_ASAP7_75t_R   g1889( .A1 (n1894), .A2 (y1110), .B (n1896), .Y (y660) );
  NOR2x1_ASAP7_75t_R   g1890( .A (n967), .B (n447), .Y (y661) );
  AND2x2_ASAP7_75t_R   g1891( .A (n443), .B (n466), .Y (y662) );
  AND2x2_ASAP7_75t_R   g1892( .A (n79), .B (n1572), .Y (n1900) );
  NOR2x1_ASAP7_75t_R   g1893( .A (n12), .B (n1900), .Y (y1134) );
  AO21x1_ASAP7_75t_R   g1894( .A1 (n12), .A2 (n1900), .B (y1134), .Y (y663) );
  NAND2x1_ASAP7_75t_R  g1895( .A (n16), .B (n1163), .Y (n1903) );
  AND2x2_ASAP7_75t_R   g1896( .A (n443), .B (n1903), .Y (y664) );
  AND2x2_ASAP7_75t_R   g1897( .A (n1115), .B (n466), .Y (y665) );
  AND3x1_ASAP7_75t_R   g1898( .A (n546), .B (y3852), .C (n466), .Y (y666) );
  AND3x1_ASAP7_75t_R   g1899( .A (y2079), .B (x4), .C (x1), .Y (n1907) );
  AO21x1_ASAP7_75t_R   g1900( .A1 (n1093), .A2 (n466), .B (n1907), .Y (y667) );
  AO21x1_ASAP7_75t_R   g1901( .A1 (n466), .A2 (x0), .B (n231), .Y (y668) );
  AO21x1_ASAP7_75t_R   g1902( .A1 (n15), .A2 (x5), .B (n143), .Y (n1910) );
  AND3x1_ASAP7_75t_R   g1903( .A (n15), .B (x1), .C (x0), .Y (n1911) );
  NAND2x1_ASAP7_75t_R  g1904( .A (x5), .B (n1911), .Y (n1912) );
  OA21x2_ASAP7_75t_R   g1905( .A1 (n1404), .A2 (n1910), .B (n1912), .Y (y669) );
  AO21x1_ASAP7_75t_R   g1906( .A1 (n466), .A2 (x0), .B (n1095), .Y (y670) );
  AO21x1_ASAP7_75t_R   g1907( .A1 (n16), .A2 (n1775), .B (n1083), .Y (y671) );
  AO21x1_ASAP7_75t_R   g1908( .A1 (n1082), .A2 (x0), .B (n1095), .Y (y673) );
  AO21x1_ASAP7_75t_R   g1909( .A1 (n12), .A2 (n22), .B (n16), .Y (n1917) );
  AO21x1_ASAP7_75t_R   g1910( .A1 (y2079), .A2 (n1917), .B (n1132), .Y (y674) );
  AO32x1_ASAP7_75t_R   g1911( .A1 (x0), .A2 (n466), .A3 (n546), .B1 (n12), .B2 (n961), .Y (y675) );
  AND2x2_ASAP7_75t_R   g1912( .A (n466), .B (n436), .Y (n1920) );
  INVx1_ASAP7_75t_R    g1913( .A (n1920), .Y (n1921) );
  AO32x1_ASAP7_75t_R   g1914( .A1 (y2079), .A2 (n1921), .A3 (n976), .B1 (n977), .B2 (n546), .Y (y676) );
  INVx1_ASAP7_75t_R    g1915( .A (n999), .Y (n1923) );
  AND3x1_ASAP7_75t_R   g1916( .A (n1923), .B (n310), .C (y2079), .Y (n1924) );
  AO21x1_ASAP7_75t_R   g1917( .A1 (n1000), .A2 (x0), .B (n1924), .Y (y677) );
  AO21x1_ASAP7_75t_R   g1918( .A1 (n1000), .A2 (x0), .B (n231), .Y (y678) );
  INVx1_ASAP7_75t_R    g1919( .A (y1281), .Y (n1927) );
  NAND2x1_ASAP7_75t_R  g1920( .A (n16), .B (n1927), .Y (n1928) );
  AND3x1_ASAP7_75t_R   g1921( .A (n1928), .B (n451), .C (n219), .Y (y679) );
  AO21x1_ASAP7_75t_R   g1922( .A1 (n1196), .A2 (x0), .B (n468), .Y (y680) );
  AND2x2_ASAP7_75t_R   g1923( .A (n1046), .B (n1047), .Y (y681) );
  AO21x1_ASAP7_75t_R   g1924( .A1 (n527), .A2 (y2079), .B (x0), .Y (n1932) );
  AND2x2_ASAP7_75t_R   g1925( .A (n1196), .B (n1932), .Y (y682) );
  AND2x2_ASAP7_75t_R   g1926( .A (n1196), .B (y1894), .Y (y939) );
  AND2x2_ASAP7_75t_R   g1927( .A (n1831), .B (y939), .Y (y683) );
  AO21x1_ASAP7_75t_R   g1928( .A1 (n437), .A2 (y2079), .B (x0), .Y (y2464) );
  AND2x2_ASAP7_75t_R   g1929( .A (y2464), .B (n1216), .Y (y684) );
  AND3x1_ASAP7_75t_R   g1930( .A (n1370), .B (n1196), .C (y1894), .Y (y685) );
  NAND2x1_ASAP7_75t_R  g1931( .A (n724), .B (y3377), .Y (n1939) );
  INVx1_ASAP7_75t_R    g1932( .A (n1939), .Y (y1445) );
  AO21x1_ASAP7_75t_R   g1933( .A1 (y1445), .A2 (n382), .B (x0), .Y (y686) );
  NAND2x1_ASAP7_75t_R  g1934( .A (n16), .B (n934), .Y (n1942) );
  AND3x1_ASAP7_75t_R   g1935( .A (n1942), .B (y1894), .C (n1370), .Y (y687) );
  AND2x2_ASAP7_75t_R   g1936( .A (n1213), .B (y1894), .Y (y688) );
  AO21x1_ASAP7_75t_R   g1937( .A1 (n1762), .A2 (n352), .B (n143), .Y (y690) );
  AO21x1_ASAP7_75t_R   g1938( .A1 (n315), .A2 (n16), .B (y2079), .Y (n1946) );
  AO21x1_ASAP7_75t_R   g1939( .A1 (x0), .A2 (x1), .B (n1946), .Y (y691) );
  AND2x2_ASAP7_75t_R   g1940( .A (n490), .B (y2079), .Y (n1948) );
  AO21x1_ASAP7_75t_R   g1941( .A1 (n1188), .A2 (n1210), .B (n1948), .Y (y692) );
  AO21x1_ASAP7_75t_R   g1942( .A1 (n12), .A2 (n22), .B (x1), .Y (n1950) );
  AO21x1_ASAP7_75t_R   g1943( .A1 (n970), .A2 (n1950), .B (n529), .Y (y693) );
  INVx1_ASAP7_75t_R    g1944( .A (n507), .Y (n1952) );
  AO21x1_ASAP7_75t_R   g1945( .A1 (n1952), .A2 (n765), .B (n989), .Y (y694) );
  OR3x1_ASAP7_75t_R    g1946( .A (x0), .B (x1), .C (x5), .Y (n1954) );
  AND2x2_ASAP7_75t_R   g1947( .A (y691), .B (n1954), .Y (y695) );
  AO21x1_ASAP7_75t_R   g1948( .A1 (n16), .A2 (n1851), .B (n1208), .Y (n1956) );
  INVx1_ASAP7_75t_R    g1949( .A (n1956), .Y (n1957) );
  AO21x1_ASAP7_75t_R   g1950( .A1 (y9), .A2 (n529), .B (n1957), .Y (y696) );
  NOR2x1_ASAP7_75t_R   g1951( .A (n227), .B (n388), .Y (n1959) );
  AND3x1_ASAP7_75t_R   g1952( .A (n315), .B (n16), .C (x5), .Y (n1960) );
  OR3x1_ASAP7_75t_R    g1953( .A (n1959), .B (n1960), .C (y863), .Y (y697) );
  OAI21x1_ASAP7_75t_R  g1954( .A1 (n58), .A2 (n507), .B (n1802), .Y (y699) );
  AO21x1_ASAP7_75t_R   g1955( .A1 (y2079), .A2 (x4), .B (n43), .Y (n1963) );
  AO21x1_ASAP7_75t_R   g1956( .A1 (x1), .A2 (n58), .B (n1963), .Y (n1964) );
  AND2x2_ASAP7_75t_R   g1957( .A (n1964), .B (n1853), .Y (y700) );
  AND2x2_ASAP7_75t_R   g1958( .A (y694), .B (n455), .Y (y701) );
  AO21x1_ASAP7_75t_R   g1959( .A1 (x0), .A2 (x1), .B (n1095), .Y (n1967) );
  AO21x1_ASAP7_75t_R   g1960( .A1 (n315), .A2 (n776), .B (n1967), .Y (y702) );
  AO21x1_ASAP7_75t_R   g1961( .A1 (n22), .A2 (y2079), .B (x1), .Y (n1969) );
  NAND2x1_ASAP7_75t_R  g1962( .A (n12), .B (n1969), .Y (n1970) );
  OR3x1_ASAP7_75t_R    g1963( .A (n315), .B (y2079), .C (x1), .Y (n1971) );
  AND2x2_ASAP7_75t_R   g1964( .A (n1970), .B (n1971), .Y (y703) );
  OA21x2_ASAP7_75t_R   g1965( .A1 (n25), .A2 (n315), .B (n219), .Y (y704) );
  OR3x1_ASAP7_75t_R    g1966( .A (n529), .B (n306), .C (x1), .Y (n1974) );
  AND2x2_ASAP7_75t_R   g1967( .A (n1974), .B (n219), .Y (y705) );
  AO21x1_ASAP7_75t_R   g1968( .A1 (n22), .A2 (n700), .B (n538), .Y (y706) );
  AO21x1_ASAP7_75t_R   g1969( .A1 (n455), .A2 (n143), .B (n231), .Y (n1977) );
  AO21x1_ASAP7_75t_R   g1970( .A1 (n315), .A2 (n776), .B (n1977), .Y (y707) );
  OR3x1_ASAP7_75t_R    g1971( .A (y3758), .B (n437), .C (x0), .Y (y708) );
  AO21x1_ASAP7_75t_R   g1972( .A1 (x1), .A2 (x4), .B (x5), .Y (n1980) );
  XOR2x2_ASAP7_75t_R   g1973( .A (n1956), .B (n1980), .Y (y709) );
  AND2x2_ASAP7_75t_R   g1974( .A (n457), .B (x0), .Y (y3047) );
  AO21x1_ASAP7_75t_R   g1975( .A1 (n419), .A2 (n43), .B (y3047), .Y (y710) );
  AND2x2_ASAP7_75t_R   g1976( .A (n1215), .B (n219), .Y (n1984) );
  AO21x1_ASAP7_75t_R   g1977( .A1 (n776), .A2 (n315), .B (n1984), .Y (y711) );
  AND2x2_ASAP7_75t_R   g1978( .A (n1971), .B (n219), .Y (y2280) );
  AND2x2_ASAP7_75t_R   g1979( .A (n1064), .B (y2280), .Y (y712) );
  AO221x2_ASAP7_75t_R  g1980( .A1 (n315), .A2 (n312), .B1 (y195), .B2 (x4), .C (y772), .Y (y713) );
  INVx1_ASAP7_75t_R    g1981( .A (n1125), .Y (n1989) );
  NOR2x1_ASAP7_75t_R   g1982( .A (n1012), .B (n1989), .Y (y714) );
  OA21x2_ASAP7_75t_R   g1983( .A1 (x0), .A2 (n552), .B (n1246), .Y (y715) );
  INVx1_ASAP7_75t_R    g1984( .A (n578), .Y (n1992) );
  OA21x2_ASAP7_75t_R   g1985( .A1 (n1992), .A2 (x0), .B (n1246), .Y (y716) );
  AO32x1_ASAP7_75t_R   g1986( .A1 (n534), .A2 (y3852), .A3 (n1851), .B1 (n315), .B2 (n312), .Y (y717) );
  AND2x2_ASAP7_75t_R   g1987( .A (n25), .B (x0), .Y (n1995) );
  AO21x1_ASAP7_75t_R   g1988( .A1 (n776), .A2 (n315), .B (n1995), .Y (y718) );
  AO21x1_ASAP7_75t_R   g1989( .A1 (x4), .A2 (x5), .B (x3), .Y (n1997) );
  OA21x2_ASAP7_75t_R   g1990( .A1 (y3758), .A2 (n84), .B (n1997), .Y (y719) );
  NOR2x1_ASAP7_75t_R   g1991( .A (n1245), .B (n1189), .Y (y720) );
  AO21x1_ASAP7_75t_R   g1992( .A1 (n1046), .A2 (x0), .B (n344), .Y (y721) );
  AND3x1_ASAP7_75t_R   g1993( .A (n527), .B (n12), .C (x5), .Y (n2001) );
  AO21x1_ASAP7_75t_R   g1994( .A1 (n497), .A2 (x0), .B (n2001), .Y (y722) );
  OR3x1_ASAP7_75t_R    g1995( .A (n529), .B (n12), .C (n544), .Y (n2003) );
  OA21x2_ASAP7_75t_R   g1996( .A1 (x0), .A2 (n552), .B (n2003), .Y (y723) );
  AND3x1_ASAP7_75t_R   g1997( .A (n856), .B (n16), .C (x0), .Y (n2005) );
  INVx1_ASAP7_75t_R    g1998( .A (n2005), .Y (n2006) );
  AND2x2_ASAP7_75t_R   g1999( .A (n2006), .B (y22), .Y (y724) );
  AO21x1_ASAP7_75t_R   g2000( .A1 (n22), .A2 (x1), .B (n12), .Y (n2008) );
  INVx1_ASAP7_75t_R    g2001( .A (n2008), .Y (n2009) );
  OA21x2_ASAP7_75t_R   g2002( .A1 (n970), .A2 (n2009), .B (n1971), .Y (y725) );
  AO21x1_ASAP7_75t_R   g2003( .A1 (y2079), .A2 (n22), .B (y863), .Y (y2659) );
  AO21x1_ASAP7_75t_R   g2004( .A1 (n606), .A2 (n12), .B (y2659), .Y (y726) );
  INVx1_ASAP7_75t_R    g2005( .A (n429), .Y (n2013) );
  AO21x1_ASAP7_75t_R   g2006( .A1 (n2013), .A2 (n16), .B (n143), .Y (y727) );
  AND3x1_ASAP7_75t_R   g2007( .A (n1246), .B (n219), .C (n1265), .Y (y728) );
  AO21x1_ASAP7_75t_R   g2008( .A1 (n388), .A2 (n28), .B (x0), .Y (n2016) );
  INVx1_ASAP7_75t_R    g2009( .A (n2016), .Y (n2017) );
  AO21x1_ASAP7_75t_R   g2010( .A1 (n2017), .A2 (n16), .B (n143), .Y (y729) );
  INVx1_ASAP7_75t_R    g2011( .A (n1817), .Y (n2019) );
  AO21x1_ASAP7_75t_R   g2012( .A1 (y3852), .A2 (n352), .B (x4), .Y (n2020) );
  AO21x1_ASAP7_75t_R   g2013( .A1 (n12), .A2 (n419), .B (y2498), .Y (n2021) );
  AO32x1_ASAP7_75t_R   g2014( .A1 (n16), .A2 (n2019), .A3 (n2020), .B1 (x1), .B2 (n2021), .Y (n2022) );
  INVx1_ASAP7_75t_R    g2015( .A (n2022), .Y (y730) );
  OR3x1_ASAP7_75t_R    g2016( .A (y2466), .B (n16), .C (n12), .Y (n2024) );
  NAND2x1_ASAP7_75t_R  g2017( .A (n510), .B (n512), .Y (n2025) );
  NAND2x1_ASAP7_75t_R  g2018( .A (n2024), .B (n2025), .Y (y731) );
  AO21x1_ASAP7_75t_R   g2019( .A1 (x0), .A2 (x4), .B (x5), .Y (n2027) );
  INVx1_ASAP7_75t_R    g2020( .A (n1950), .Y (n2028) );
  OA222x2_ASAP7_75t_R  g2021( .A1 (n2027), .A2 (n2028), .B1 (x0), .B2 (n16), .C1 (n457), .C2 (n2013), .Y (y732) );
  AO21x1_ASAP7_75t_R   g2022( .A1 (n419), .A2 (n143), .B (n929), .Y (y733) );
  NAND2x1_ASAP7_75t_R  g2023( .A (n16), .B (n429), .Y (n2031) );
  AND3x1_ASAP7_75t_R   g2024( .A (n2031), .B (n219), .C (n419), .Y (y734) );
  AO21x1_ASAP7_75t_R   g2025( .A1 (n175), .A2 (y2079), .B (y863), .Y (y735) );
  NAND2x1_ASAP7_75t_R  g2026( .A (n180), .B (n740), .Y (y736) );
  AND2x2_ASAP7_75t_R   g2027( .A (n1235), .B (y2813), .Y (y737) );
  NOR2x1_ASAP7_75t_R   g2028( .A (n12), .B (n1190), .Y (n2036) );
  AO21x1_ASAP7_75t_R   g2029( .A1 (n998), .A2 (n12), .B (n2036), .Y (y738) );
  AO21x1_ASAP7_75t_R   g2030( .A1 (n16), .A2 (x0), .B (x2), .Y (n2038) );
  AO21x1_ASAP7_75t_R   g2031( .A1 (n2038), .A2 (y2079), .B (n1778), .Y (y739) );
  OR3x1_ASAP7_75t_R    g2032( .A (n43), .B (x5), .C (x2), .Y (n2040) );
  AND2x2_ASAP7_75t_R   g2033( .A (n2040), .B (n1782), .Y (y740) );
  AND2x2_ASAP7_75t_R   g2034( .A (n707), .B (n994), .Y (y742) );
  AND2x2_ASAP7_75t_R   g2035( .A (y1283), .B (n187), .Y (y743) );
  AO21x1_ASAP7_75t_R   g2036( .A1 (n1269), .A2 (y9), .B (n143), .Y (y744) );
  AND2x2_ASAP7_75t_R   g2037( .A (n1383), .B (n1340), .Y (y745) );
  AND3x1_ASAP7_75t_R   g2038( .A (n1340), .B (y195), .C (n497), .Y (y746) );
  AND3x1_ASAP7_75t_R   g2039( .A (n363), .B (n15), .C (n16), .Y (n2047) );
  AO21x1_ASAP7_75t_R   g2040( .A1 (y741), .A2 (n1265), .B (n2047), .Y (y747) );
  AO21x1_ASAP7_75t_R   g2041( .A1 (n360), .A2 (n290), .B (y2079), .Y (n2049) );
  INVx1_ASAP7_75t_R    g2042( .A (n2049), .Y (n2050) );
  AND3x1_ASAP7_75t_R   g2043( .A (n360), .B (n290), .C (y2079), .Y (n2051) );
  OR3x1_ASAP7_75t_R    g2044( .A (n2050), .B (n2051), .C (x0), .Y (y748) );
  AO21x1_ASAP7_75t_R   g2045( .A1 (n1269), .A2 (y9), .B (n1778), .Y (y749) );
  INVx1_ASAP7_75t_R    g2046( .A (n1980), .Y (n2054) );
  AO21x1_ASAP7_75t_R   g2047( .A1 (x0), .A2 (x1), .B (n2054), .Y (y750) );
  AO21x1_ASAP7_75t_R   g2048( .A1 (x0), .A2 (x1), .B (n1924), .Y (y751) );
  AND2x2_ASAP7_75t_R   g2049( .A (n497), .B (n1424), .Y (y752) );
  AND2x2_ASAP7_75t_R   g2050( .A (n1125), .B (n604), .Y (y753) );
  AO21x1_ASAP7_75t_R   g2051( .A1 (n15), .A2 (x0), .B (x5), .Y (n2059) );
  INVx1_ASAP7_75t_R    g2052( .A (n2059), .Y (n2060) );
  AO21x1_ASAP7_75t_R   g2053( .A1 (n2060), .A2 (n16), .B (n143), .Y (y754) );
  AND2x2_ASAP7_75t_R   g2054( .A (n496), .B (n1218), .Y (y755) );
  AO21x1_ASAP7_75t_R   g2055( .A1 (y2079), .A2 (x4), .B (n12), .Y (n2063) );
  NAND2x1_ASAP7_75t_R  g2056( .A (n2063), .B (n312), .Y (y756) );
  AO21x1_ASAP7_75t_R   g2057( .A1 (x0), .A2 (x1), .B (n705), .Y (y757) );
  AO21x1_ASAP7_75t_R   g2058( .A1 (y2079), .A2 (n1426), .B (n1292), .Y (y758) );
  NOR2x1_ASAP7_75t_R   g2059( .A (x5), .B (n241), .Y (n2067) );
  NAND2x1_ASAP7_75t_R  g2060( .A (x1), .B (n692), .Y (n2068) );
  OR3x1_ASAP7_75t_R    g2061( .A (x0), .B (x2), .C (x5), .Y (n2069) );
  INVx1_ASAP7_75t_R    g2062( .A (n2069), .Y (n2070) );
  OA22x2_ASAP7_75t_R   g2063( .A1 (x1), .A2 (n2067), .B1 (n2068), .B2 (n2070), .Y (y759) );
  AO21x1_ASAP7_75t_R   g2064( .A1 (y2079), .A2 (n52), .B (n761), .Y (n2072) );
  AND2x2_ASAP7_75t_R   g2065( .A (n2072), .B (n14), .Y (n2073) );
  NOR2x1_ASAP7_75t_R   g2066( .A (n481), .B (n2073), .Y (y760) );
  AND3x1_ASAP7_75t_R   g2067( .A (n714), .B (n1438), .C (n497), .Y (y761) );
  AO21x1_ASAP7_75t_R   g2068( .A1 (n1265), .A2 (n143), .B (n231), .Y (y762) );
  OA21x2_ASAP7_75t_R   g2069( .A1 (x1), .A2 (n2067), .B (n2068), .Y (y763) );
  AO21x1_ASAP7_75t_R   g2070( .A1 (n16), .A2 (y2079), .B (n143), .Y (y1356) );
  AND2x2_ASAP7_75t_R   g2071( .A (n714), .B (y1356), .Y (y764) );
  AND2x2_ASAP7_75t_R   g2072( .A (n665), .B (n219), .Y (y765) );
  AO21x1_ASAP7_75t_R   g2073( .A1 (n497), .A2 (x0), .B (y2466), .Y (y766) );
  AND2x2_ASAP7_75t_R   g2074( .A (n1047), .B (n994), .Y (y767) );
  AO21x1_ASAP7_75t_R   g2075( .A1 (n25), .A2 (x0), .B (n344), .Y (y768) );
  AND2x2_ASAP7_75t_R   g2076( .A (n1047), .B (n25), .Y (y769) );
  AO21x1_ASAP7_75t_R   g2077( .A1 (n1210), .A2 (n1188), .B (n529), .Y (n2085) );
  AO21x1_ASAP7_75t_R   g2078( .A1 (n1956), .A2 (y2079), .B (n2085), .Y (y770) );
  AND2x2_ASAP7_75t_R   g2079( .A (n497), .B (n1188), .Y (y771) );
  AO21x1_ASAP7_75t_R   g2080( .A1 (n665), .A2 (x0), .B (n2070), .Y (y774) );
  AO21x1_ASAP7_75t_R   g2081( .A1 (n665), .A2 (x0), .B (n1315), .Y (y775) );
  INVx1_ASAP7_75t_R    g2082( .A (n743), .Y (n2090) );
  AO21x1_ASAP7_75t_R   g2083( .A1 (n665), .A2 (x0), .B (n2090), .Y (y776) );
  OR3x1_ASAP7_75t_R    g2084( .A (n993), .B (n12), .C (n1339), .Y (n2092) );
  INVx1_ASAP7_75t_R    g2085( .A (n2092), .Y (y777) );
  AND3x1_ASAP7_75t_R   g2086( .A (n714), .B (n497), .C (n1457), .Y (y778) );
  AO21x1_ASAP7_75t_R   g2087( .A1 (n15), .A2 (y2079), .B (x1), .Y (n2095) );
  AND2x2_ASAP7_75t_R   g2088( .A (n2095), .B (x0), .Y (n2096) );
  INVx1_ASAP7_75t_R    g2089( .A (n1324), .Y (n2097) );
  AO21x1_ASAP7_75t_R   g2090( .A1 (n1340), .A2 (n2096), .B (n2097), .Y (y779) );
  INVx1_ASAP7_75t_R    g2091( .A (n1385), .Y (n2099) );
  AO21x1_ASAP7_75t_R   g2092( .A1 (n1265), .A2 (y863), .B (n2099), .Y (y780) );
  NAND2x1_ASAP7_75t_R  g2093( .A (n492), .B (n490), .Y (y781) );
  AO21x1_ASAP7_75t_R   g2094( .A1 (n363), .A2 (n16), .B (n143), .Y (y873) );
  AND2x2_ASAP7_75t_R   g2095( .A (y873), .B (n1265), .Y (y782) );
  OR3x1_ASAP7_75t_R    g2096( .A (n347), .B (y2079), .C (x0), .Y (n2104) );
  AND2x2_ASAP7_75t_R   g2097( .A (n1161), .B (n2104), .Y (y783) );
  AO21x1_ASAP7_75t_R   g2098( .A1 (n1265), .A2 (n143), .B (n1060), .Y (y784) );
  INVx1_ASAP7_75t_R    g2099( .A (n947), .Y (n2107) );
  AO21x1_ASAP7_75t_R   g2100( .A1 (n2107), .A2 (y2079), .B (y863), .Y (y785) );
  AO21x1_ASAP7_75t_R   g2101( .A1 (n546), .A2 (y3127), .B (n1155), .Y (y786) );
  NAND2x1_ASAP7_75t_R  g2102( .A (n1358), .B (n1356), .Y (y787) );
  AND2x2_ASAP7_75t_R   g2103( .A (y787), .B (n228), .Y (y788) );
  AO21x1_ASAP7_75t_R   g2104( .A1 (n1572), .A2 (n143), .B (n1874), .Y (y789) );
  INVx1_ASAP7_75t_R    g2105( .A (n674), .Y (n2113) );
  OA21x2_ASAP7_75t_R   g2106( .A1 (n2113), .A2 (n1874), .B (x0), .Y (y790) );
  AO21x1_ASAP7_75t_R   g2107( .A1 (n64), .A2 (n1546), .B (x0), .Y (y791) );
  INVx1_ASAP7_75t_R    g2108( .A (n1911), .Y (n2116) );
  AO21x1_ASAP7_75t_R   g2109( .A1 (x0), .A2 (x1), .B (n15), .Y (n2117) );
  AO21x1_ASAP7_75t_R   g2110( .A1 (n2116), .A2 (n2117), .B (y2079), .Y (y792) );
  AND2x2_ASAP7_75t_R   g2111( .A (y2813), .B (x2), .Y (n2119) );
  OR3x1_ASAP7_75t_R    g2112( .A (n1541), .B (y2093), .C (n2119), .Y (y793) );
  AO21x1_ASAP7_75t_R   g2113( .A1 (x1), .A2 (n276), .B (n1454), .Y (n2121) );
  AND3x1_ASAP7_75t_R   g2114( .A (n12), .B (n15), .C (x1), .Y (n2122) );
  INVx1_ASAP7_75t_R    g2115( .A (n2122), .Y (n2123) );
  AO22x1_ASAP7_75t_R   g2116( .A1 (x5), .A2 (n2121), .B1 (y2079), .B2 (n2123), .Y (y794) );
  OR3x1_ASAP7_75t_R    g2117( .A (n143), .B (y2079), .C (x2), .Y (n2125) );
  INVx1_ASAP7_75t_R    g2118( .A (n2125), .Y (n2126) );
  AO21x1_ASAP7_75t_R   g2119( .A1 (n1502), .A2 (n1782), .B (n2126), .Y (y795) );
  OR3x1_ASAP7_75t_R    g2120( .A (y863), .B (y2079), .C (n15), .Y (n2128) );
  AND2x2_ASAP7_75t_R   g2121( .A (n1232), .B (n2128), .Y (y796) );
  AO32x1_ASAP7_75t_R   g2122( .A1 (n173), .A2 (n1385), .A3 (n15), .B1 (x2), .B2 (y2813), .Y (y797) );
  OR3x1_ASAP7_75t_R    g2123( .A (n227), .B (y2079), .C (n22), .Y (n2131) );
  AO21x1_ASAP7_75t_R   g2124( .A1 (n1310), .A2 (n2131), .B (y863), .Y (y798) );
  AO21x1_ASAP7_75t_R   g2125( .A1 (x5), .A2 (n12), .B (n63), .Y (n2133) );
  OR3x1_ASAP7_75t_R    g2126( .A (n143), .B (y2079), .C (n15), .Y (n2134) );
  AND2x2_ASAP7_75t_R   g2127( .A (n2133), .B (n2134), .Y (y799) );
  AO21x1_ASAP7_75t_R   g2128( .A1 (n12), .A2 (y2079), .B (x2), .Y (n2136) );
  INVx1_ASAP7_75t_R    g2129( .A (n2136), .Y (n2137) );
  AO21x1_ASAP7_75t_R   g2130( .A1 (n2137), .A2 (n144), .B (n1269), .Y (n2138) );
  AO21x1_ASAP7_75t_R   g2131( .A1 (x2), .A2 (n1819), .B (n2138), .Y (y800) );
  AO21x1_ASAP7_75t_R   g2132( .A1 (n12), .A2 (x5), .B (x2), .Y (n2140) );
  AO21x1_ASAP7_75t_R   g2133( .A1 (n352), .A2 (n16), .B (n2140), .Y (n2141) );
  AND2x2_ASAP7_75t_R   g2134( .A (n2141), .B (n2134), .Y (y801) );
  AO21x1_ASAP7_75t_R   g2135( .A1 (n173), .A2 (n1646), .B (n2119), .Y (y802) );
  OA21x2_ASAP7_75t_R   g2136( .A1 (y741), .A2 (n1646), .B (n1912), .Y (y803) );
  NAND2x1_ASAP7_75t_R  g2137( .A (n15), .B (n988), .Y (n2145) );
  INVx1_ASAP7_75t_R    g2138( .A (n2145), .Y (n2146) );
  NOR2x1_ASAP7_75t_R   g2139( .A (n15), .B (n988), .Y (n2147) );
  OR3x1_ASAP7_75t_R    g2140( .A (n2146), .B (n2147), .C (y2196), .Y (y804) );
  OR3x1_ASAP7_75t_R    g2141( .A (n2126), .B (n2147), .C (y2196), .Y (y805) );
  AO21x1_ASAP7_75t_R   g2142( .A1 (y3852), .A2 (x1), .B (n835), .Y (n2150) );
  AND2x2_ASAP7_75t_R   g2143( .A (n2150), .B (n2116), .Y (y806) );
  AO32x1_ASAP7_75t_R   g2144( .A1 (n757), .A2 (n173), .A3 (n1385), .B1 (n103), .B2 (x0), .Y (y807) );
  AND2x2_ASAP7_75t_R   g2145( .A (n2150), .B (n2133), .Y (y808) );
  NAND2x1_ASAP7_75t_R  g2146( .A (n97), .B (n352), .Y (n2154) );
  AO21x1_ASAP7_75t_R   g2147( .A1 (n2154), .A2 (n988), .B (n2147), .Y (y809) );
  AND3x1_ASAP7_75t_R   g2148( .A (y3852), .B (n994), .C (x2), .Y (n2156) );
  AO21x1_ASAP7_75t_R   g2149( .A1 (n1106), .A2 (n1454), .B (n2156), .Y (y810) );
  AO21x1_ASAP7_75t_R   g2150( .A1 (x0), .A2 (x2), .B (n16), .Y (n2158) );
  AO21x1_ASAP7_75t_R   g2151( .A1 (n64), .A2 (n2158), .B (n1565), .Y (y811) );
  NOR2x1_ASAP7_75t_R   g2152( .A (n12), .B (n99), .Y (n2160) );
  OR3x1_ASAP7_75t_R    g2153( .A (n771), .B (n2160), .C (n241), .Y (y812) );
  INVx1_ASAP7_75t_R    g2154( .A (n1778), .Y (n2162) );
  AO21x1_ASAP7_75t_R   g2155( .A1 (n16), .A2 (y2079), .B (x2), .Y (n2163) );
  INVx1_ASAP7_75t_R    g2156( .A (n2163), .Y (n2164) );
  AND2x2_ASAP7_75t_R   g2157( .A (y1356), .B (x2), .Y (n2165) );
  AO21x1_ASAP7_75t_R   g2158( .A1 (n2162), .A2 (n2164), .B (n2165), .Y (y813) );
  OA21x2_ASAP7_75t_R   g2159( .A1 (y757), .A2 (n1646), .B (n1912), .Y (y814) );
  OA21x2_ASAP7_75t_R   g2160( .A1 (n15), .A2 (y1356), .B (n2116), .Y (y815) );
  AND3x1_ASAP7_75t_R   g2161( .A (x0), .B (x1), .C (x2), .Y (n2169) );
  OR3x1_ASAP7_75t_R    g2162( .A (n2126), .B (n2169), .C (n231), .Y (y816) );
  AO21x1_ASAP7_75t_R   g2163( .A1 (n144), .A2 (n2137), .B (n2165), .Y (y817) );
  AO21x1_ASAP7_75t_R   g2164( .A1 (x1), .A2 (x2), .B (y2079), .Y (n2172) );
  AND2x2_ASAP7_75t_R   g2165( .A (n2172), .B (x0), .Y (n2173) );
  AO21x1_ASAP7_75t_R   g2166( .A1 (n15), .A2 (n180), .B (n2173), .Y (y818) );
  AO21x1_ASAP7_75t_R   g2167( .A1 (n12), .A2 (n72), .B (n1549), .Y (n2175) );
  AO32x1_ASAP7_75t_R   g2168( .A1 (n16), .A2 (n1550), .A3 (n1484), .B1 (n1482), .B2 (n2175), .Y (n2176) );
  INVx1_ASAP7_75t_R    g2169( .A (n2176), .Y (y819) );
  AND3x1_ASAP7_75t_R   g2170( .A (n700), .B (n144), .C (n15), .Y (n2178) );
  AO21x1_ASAP7_75t_R   g2171( .A1 (n2172), .A2 (x0), .B (n2178), .Y (y820) );
  AO21x1_ASAP7_75t_R   g2172( .A1 (x0), .A2 (x5), .B (n16), .Y (n2180) );
  INVx1_ASAP7_75t_R    g2173( .A (n2180), .Y (n2181) );
  NAND2x1_ASAP7_75t_R  g2174( .A (x2), .B (n180), .Y (n2182) );
  OA21x2_ASAP7_75t_R   g2175( .A1 (n2181), .A2 (n750), .B (n2182), .Y (y821) );
  AO21x1_ASAP7_75t_R   g2176( .A1 (y2079), .A2 (n290), .B (n297), .Y (n2184) );
  OR3x1_ASAP7_75t_R    g2177( .A (n2184), .B (n1158), .C (x0), .Y (y822) );
  OA21x2_ASAP7_75t_R   g2178( .A1 (n993), .A2 (n707), .B (n1246), .Y (y823) );
  AO21x1_ASAP7_75t_R   g2179( .A1 (n2172), .A2 (x0), .B (n128), .Y (y1625) );
  AO21x1_ASAP7_75t_R   g2180( .A1 (n481), .A2 (n15), .B (y1625), .Y (y824) );
  AO21x1_ASAP7_75t_R   g2181( .A1 (y2079), .A2 (x2), .B (n16), .Y (n2189) );
  NOR2x1_ASAP7_75t_R   g2182( .A (x0), .B (n2189), .Y (n2190) );
  NOR2x1_ASAP7_75t_R   g2183( .A (n1245), .B (n2190), .Y (y825) );
  AO21x1_ASAP7_75t_R   g2184( .A1 (n144), .A2 (n1646), .B (n2173), .Y (y826) );
  AND3x1_ASAP7_75t_R   g2185( .A (n97), .B (n1336), .C (x0), .Y (n2193) );
  AO21x1_ASAP7_75t_R   g2186( .A1 (n1106), .A2 (n1454), .B (n2193), .Y (y827) );
  OR3x1_ASAP7_75t_R    g2187( .A (n856), .B (n12), .C (n16), .Y (n2195) );
  NAND2x1_ASAP7_75t_R  g2188( .A (n2195), .B (n1598), .Y (y828) );
  AO21x1_ASAP7_75t_R   g2189( .A1 (n497), .A2 (n276), .B (n1454), .Y (y829) );
  AO21x1_ASAP7_75t_R   g2190( .A1 (n2163), .A2 (y772), .B (n2178), .Y (y830) );
  AO21x1_ASAP7_75t_R   g2191( .A1 (x5), .A2 (n16), .B (n1469), .Y (n2199) );
  NAND2x1_ASAP7_75t_R  g2192( .A (n2199), .B (n2145), .Y (y831) );
  AND3x1_ASAP7_75t_R   g2193( .A (n2116), .B (n2134), .C (n583), .Y (y832) );
  AND2x2_ASAP7_75t_R   g2194( .A (n1106), .B (n1454), .Y (n2202) );
  AO21x1_ASAP7_75t_R   g2195( .A1 (n497), .A2 (n276), .B (n2202), .Y (y833) );
  OR3x1_ASAP7_75t_R    g2196( .A (n590), .B (n22), .C (n58), .Y (n2204) );
  AND2x2_ASAP7_75t_R   g2197( .A (n2204), .B (n980), .Y (y834) );
  AO21x1_ASAP7_75t_R   g2198( .A1 (n497), .A2 (n276), .B (n2126), .Y (y835) );
  AO32x1_ASAP7_75t_R   g2199( .A1 (n1954), .A2 (n1291), .A3 (n15), .B1 (x2), .B2 (y873), .Y (y836) );
  AO21x1_ASAP7_75t_R   g2200( .A1 (n12), .A2 (y2079), .B (n15), .Y (n2208) );
  AO21x1_ASAP7_75t_R   g2201( .A1 (n2208), .A2 (n988), .B (n2160), .Y (y837) );
  INVx1_ASAP7_75t_R    g2202( .A (n1492), .Y (n2210) );
  AO21x1_ASAP7_75t_R   g2203( .A1 (x0), .A2 (n16), .B (n97), .Y (n2211) );
  INVx1_ASAP7_75t_R    g2204( .A (n2211), .Y (n2212) );
  AO21x1_ASAP7_75t_R   g2205( .A1 (n16), .A2 (n2210), .B (n2212), .Y (n2213) );
  XOR2x2_ASAP7_75t_R   g2206( .A (n2213), .B (x0), .Y (y838) );
  AND3x1_ASAP7_75t_R   g2207( .A (n674), .B (n1873), .C (n12), .Y (n2215) );
  INVx1_ASAP7_75t_R    g2208( .A (n2215), .Y (y839) );
  NAND2x1_ASAP7_75t_R  g2209( .A (x1), .B (n168), .Y (n2217) );
  OR3x1_ASAP7_75t_R    g2210( .A (n81), .B (n12), .C (x1), .Y (n2218) );
  AND2x2_ASAP7_75t_R   g2211( .A (n2217), .B (n2218), .Y (y840) );
  OA21x2_ASAP7_75t_R   g2212( .A1 (n1646), .A2 (y873), .B (n1912), .Y (y841) );
  AND3x1_ASAP7_75t_R   g2213( .A (n90), .B (n17), .C (n15), .Y (n2221) );
  INVx1_ASAP7_75t_R    g2214( .A (n2221), .Y (n2222) );
  OR3x1_ASAP7_75t_R    g2215( .A (n45), .B (n12), .C (x1), .Y (n2223) );
  AND2x2_ASAP7_75t_R   g2216( .A (n2223), .B (n219), .Y (n2224) );
  AND2x2_ASAP7_75t_R   g2217( .A (n2222), .B (n2224), .Y (y842) );
  AO21x1_ASAP7_75t_R   g2218( .A1 (n15), .A2 (x5), .B (n701), .Y (n2226) );
  AO33x2_ASAP7_75t_R   g2219( .A1 (n97), .A2 (n144), .A3 (n1387), .B1 (n707), .B2 (n2226), .B3 (x1), .Y (n2227) );
  INVx1_ASAP7_75t_R    g2220( .A (n2227), .Y (y843) );
  INVx1_ASAP7_75t_R    g2221( .A (n554), .Y (n2229) );
  AO21x1_ASAP7_75t_R   g2222( .A1 (n388), .A2 (n538), .B (n2229), .Y (y844) );
  AND3x1_ASAP7_75t_R   g2223( .A (n622), .B (n64), .C (n610), .Y (n2231) );
  INVx1_ASAP7_75t_R    g2224( .A (n2223), .Y (n2232) );
  NOR2x1_ASAP7_75t_R   g2225( .A (n2231), .B (n2232), .Y (y845) );
  AO32x1_ASAP7_75t_R   g2226( .A1 (n144), .A2 (n1954), .A3 (n15), .B1 (x2), .B2 (y873), .Y (y846) );
  AO21x1_ASAP7_75t_R   g2227( .A1 (y2079), .A2 (x4), .B (n1380), .Y (n2235) );
  AO21x1_ASAP7_75t_R   g2228( .A1 (n527), .A2 (n12), .B (n2235), .Y (y847) );
  AO21x1_ASAP7_75t_R   g2229( .A1 (n583), .A2 (n746), .B (n16), .Y (n2237) );
  OA21x2_ASAP7_75t_R   g2230( .A1 (n989), .A2 (n2208), .B (n2237), .Y (y848) );
  NAND2x1_ASAP7_75t_R  g2231( .A (n15), .B (n1782), .Y (n2239) );
  OA21x2_ASAP7_75t_R   g2232( .A1 (n15), .A2 (y873), .B (n2239), .Y (y849) );
  AO21x1_ASAP7_75t_R   g2233( .A1 (n15), .A2 (x5), .B (y863), .Y (n2241) );
  AO21x1_ASAP7_75t_R   g2234( .A1 (n15), .A2 (n228), .B (n2241), .Y (n2242) );
  NAND2x1_ASAP7_75t_R  g2235( .A (x5), .B (n1231), .Y (n2243) );
  AND2x2_ASAP7_75t_R   g2236( .A (n2242), .B (n2243), .Y (y850) );
  AO21x1_ASAP7_75t_R   g2237( .A1 (n17), .A2 (x0), .B (n518), .Y (n2245) );
  INVx1_ASAP7_75t_R    g2238( .A (n2245), .Y (n2246) );
  AO21x1_ASAP7_75t_R   g2239( .A1 (n396), .A2 (n84), .B (n2246), .Y (y851) );
  AND3x1_ASAP7_75t_R   g2240( .A (n1912), .B (n2117), .C (n583), .Y (y852) );
  OA21x2_ASAP7_75t_R   g2241( .A1 (n529), .A2 (n962), .B (x0), .Y (n2249) );
  AO21x1_ASAP7_75t_R   g2242( .A1 (n12), .A2 (n1173), .B (n2249), .Y (y853) );
  AO21x1_ASAP7_75t_R   g2243( .A1 (n1242), .A2 (n271), .B (y2163), .Y (y854) );
  AO21x1_ASAP7_75t_R   g2244( .A1 (n173), .A2 (x2), .B (n1231), .Y (n2252) );
  INVx1_ASAP7_75t_R    g2245( .A (n2252), .Y (y855) );
  AO21x1_ASAP7_75t_R   g2246( .A1 (x3), .A2 (n12), .B (n63), .Y (n2254) );
  AND2x2_ASAP7_75t_R   g2247( .A (n2254), .B (n2117), .Y (y856) );
  AO21x1_ASAP7_75t_R   g2248( .A1 (n16), .A2 (n12), .B (x3), .Y (n2256) );
  AO21x1_ASAP7_75t_R   g2249( .A1 (n2256), .A2 (n271), .B (n262), .Y (y857) );
  INVx1_ASAP7_75t_R    g2250( .A (n262), .Y (n2258) );
  AO21x1_ASAP7_75t_R   g2251( .A1 (n2258), .A2 (n17), .B (n271), .Y (n2259) );
  AO21x1_ASAP7_75t_R   g2252( .A1 (x2), .A2 (n1682), .B (n2259), .Y (y858) );
  AO21x1_ASAP7_75t_R   g2253( .A1 (n137), .A2 (n72), .B (n12), .Y (n2261) );
  NOR2x1_ASAP7_75t_R   g2254( .A (n16), .B (n2261), .Y (n2262) );
  INVx1_ASAP7_75t_R    g2255( .A (n2262), .Y (n2263) );
  INVx1_ASAP7_75t_R    g2256( .A (n1391), .Y (n2264) );
  OR3x1_ASAP7_75t_R    g2257( .A (n218), .B (n2264), .C (y863), .Y (n2265) );
  AND2x2_ASAP7_75t_R   g2258( .A (n2263), .B (n2265), .Y (y859) );
  AO21x1_ASAP7_75t_R   g2259( .A1 (n665), .A2 (x0), .B (n43), .Y (y860) );
  AO32x1_ASAP7_75t_R   g2260( .A1 (n17), .A2 (n2258), .A3 (n1594), .B1 (x3), .B2 (n272), .Y (y861) );
  INVx1_ASAP7_75t_R    g2261( .A (n1237), .Y (n2269) );
  AND2x2_ASAP7_75t_R   g2262( .A (n2269), .B (y408), .Y (y862) );
  OR3x1_ASAP7_75t_R    g2263( .A (n163), .B (n164), .C (y863), .Y (n2271) );
  AND2x2_ASAP7_75t_R   g2264( .A (n2263), .B (n2271), .Y (y864) );
  OR3x1_ASAP7_75t_R    g2265( .A (n76), .B (n12), .C (n16), .Y (n2273) );
  OR3x1_ASAP7_75t_R    g2266( .A (y863), .B (n15), .C (n17), .Y (n2274) );
  AND2x2_ASAP7_75t_R   g2267( .A (n2273), .B (n2274), .Y (y865) );
  AO21x1_ASAP7_75t_R   g2268( .A1 (n17), .A2 (n15), .B (x0), .Y (n2276) );
  AO21x1_ASAP7_75t_R   g2269( .A1 (n12), .A2 (n15), .B (x3), .Y (n2277) );
  AND2x2_ASAP7_75t_R   g2270( .A (n72), .B (n2277), .Y (n2278) );
  INVx1_ASAP7_75t_R    g2271( .A (n2278), .Y (n2279) );
  NAND2x1_ASAP7_75t_R  g2272( .A (x1), .B (n2276), .Y (n2280) );
  AO32x1_ASAP7_75t_R   g2273( .A1 (x1), .A2 (n2276), .A3 (n2278), .B1 (n2279), .B2 (n2280), .Y (y866) );
  AO21x1_ASAP7_75t_R   g2274( .A1 (n1608), .A2 (n228), .B (x2), .Y (n2282) );
  AND2x2_ASAP7_75t_R   g2275( .A (n2282), .B (n2128), .Y (y867) );
  AND2x2_ASAP7_75t_R   g2276( .A (n1096), .B (y250), .Y (y868) );
  NAND2x1_ASAP7_75t_R  g2277( .A (n16), .B (n2027), .Y (n2285) );
  AND2x2_ASAP7_75t_R   g2278( .A (n2285), .B (n1970), .Y (y869) );
  NOR2x1_ASAP7_75t_R   g2279( .A (n12), .B (n544), .Y (n2287) );
  AO21x1_ASAP7_75t_R   g2280( .A1 (n12), .A2 (n544), .B (n2287), .Y (n2288) );
  OA21x2_ASAP7_75t_R   g2281( .A1 (n2288), .A2 (x2), .B (n2134), .Y (y870) );
  AO21x1_ASAP7_75t_R   g2282( .A1 (n701), .A2 (n16), .B (y863), .Y (y871) );
  OR3x1_ASAP7_75t_R    g2283( .A (n227), .B (y2079), .C (x2), .Y (n2291) );
  AND2x2_ASAP7_75t_R   g2284( .A (n221), .B (n1646), .Y (n2292) );
  AO21x1_ASAP7_75t_R   g2285( .A1 (y1283), .A2 (n2291), .B (n2292), .Y (y872) );
  AND2x2_ASAP7_75t_R   g2286( .A (n1466), .B (x1), .Y (n2294) );
  OA21x2_ASAP7_75t_R   g2287( .A1 (n773), .A2 (n2294), .B (n1912), .Y (y874) );
  AO21x1_ASAP7_75t_R   g2288( .A1 (n244), .A2 (x1), .B (n1889), .Y (n2296) );
  AND2x2_ASAP7_75t_R   g2289( .A (n2296), .B (n2116), .Y (y875) );
  INVx1_ASAP7_75t_R    g2290( .A (n1234), .Y (n2298) );
  AND2x2_ASAP7_75t_R   g2291( .A (n2298), .B (n2128), .Y (y876) );
  AND2x2_ASAP7_75t_R   g2292( .A (n2296), .B (n2133), .Y (y877) );
  OA21x2_ASAP7_75t_R   g2293( .A1 (x0), .A2 (n552), .B (n1283), .Y (y878) );
  AND2x2_ASAP7_75t_R   g2294( .A (n1782), .B (x2), .Y (n2302) );
  AO21x1_ASAP7_75t_R   g2295( .A1 (n988), .A2 (n1636), .B (n2302), .Y (y879) );
  AND2x2_ASAP7_75t_R   g2296( .A (n2296), .B (n2141), .Y (y880) );
  AO21x1_ASAP7_75t_R   g2297( .A1 (n221), .A2 (n1646), .B (n2119), .Y (y881) );
  AO21x1_ASAP7_75t_R   g2298( .A1 (n63), .A2 (x0), .B (n2122), .Y (n2306) );
  AO21x1_ASAP7_75t_R   g2299( .A1 (x0), .A2 (y2079), .B (n64), .Y (n2307) );
  OA21x2_ASAP7_75t_R   g2300( .A1 (n2306), .A2 (y2079), .B (n2307), .Y (y882) );
  NAND2x1_ASAP7_75t_R  g2301( .A (x5), .B (n185), .Y (n2309) );
  AO21x1_ASAP7_75t_R   g2302( .A1 (n2309), .A2 (n228), .B (n262), .Y (y883) );
  AND3x1_ASAP7_75t_R   g2303( .A (n12), .B (x2), .C (x5), .Y (n2311) );
  INVx1_ASAP7_75t_R    g2304( .A (n2311), .Y (n2312) );
  AO331x2_ASAP7_75t_R  g2305( .A1 (n16), .A2 (y3852), .A3 (n15), .B1 (n2140), .B2 (x1), .B3 (n2312), .C (y2196), .Y (y884) );
  OA21x2_ASAP7_75t_R   g2306( .A1 (n2288), .A2 (n103), .B (n2134), .Y (y885) );
  INVx1_ASAP7_75t_R    g2307( .A (n610), .Y (n2315) );
  OA21x2_ASAP7_75t_R   g2308( .A1 (n1208), .A2 (n2315), .B (n2134), .Y (y886) );
  INVx1_ASAP7_75t_R    g2309( .A (n488), .Y (n2317) );
  AO32x1_ASAP7_75t_R   g2310( .A1 (n2140), .A2 (n2312), .A3 (n994), .B1 (n15), .B2 (n2317), .Y (y887) );
  AO21x1_ASAP7_75t_R   g2311( .A1 (y9), .A2 (n757), .B (n143), .Y (n2319) );
  AND2x2_ASAP7_75t_R   g2312( .A (n2319), .B (n2133), .Y (y888) );
  INVx1_ASAP7_75t_R    g2313( .A (n1889), .Y (n2321) );
  NAND2x1_ASAP7_75t_R  g2314( .A (n16), .B (n2321), .Y (n2322) );
  INVx1_ASAP7_75t_R    g2315( .A (n772), .Y (n2323) );
  AO21x1_ASAP7_75t_R   g2316( .A1 (n2323), .A2 (n244), .B (n16), .Y (n2324) );
  AND2x2_ASAP7_75t_R   g2317( .A (n2322), .B (n2324), .Y (y889) );
  INVx1_ASAP7_75t_R    g2318( .A (n83), .Y (n2326) );
  AO21x1_ASAP7_75t_R   g2319( .A1 (n12), .A2 (n15), .B (y2079), .Y (n2327) );
  AO21x1_ASAP7_75t_R   g2320( .A1 (x2), .A2 (n16), .B (n610), .Y (n2328) );
  INVx1_ASAP7_75t_R    g2321( .A (n2328), .Y (n2329) );
  AO21x1_ASAP7_75t_R   g2322( .A1 (n2326), .A2 (n2327), .B (n2329), .Y (y891) );
  OR3x1_ASAP7_75t_R    g2323( .A (n2060), .B (n772), .C (x1), .Y (n2331) );
  AND2x2_ASAP7_75t_R   g2324( .A (n2331), .B (n2324), .Y (y892) );
  OA21x2_ASAP7_75t_R   g2325( .A1 (x1), .A2 (n773), .B (n2324), .Y (y893) );
  AO21x1_ASAP7_75t_R   g2326( .A1 (n23), .A2 (n513), .B (n549), .Y (y894) );
  XNOR2x2_ASAP7_75t_R  g2327( .A (n1424), .B (n1614), .Y (y895) );
  NAND2x1_ASAP7_75t_R  g2328( .A (n99), .B (n497), .Y (n2336) );
  XOR2x2_ASAP7_75t_R   g2329( .A (n2336), .B (n1536), .Y (y896) );
  AO21x1_ASAP7_75t_R   g2330( .A1 (n2323), .A2 (n1466), .B (n16), .Y (n2338) );
  OA21x2_ASAP7_75t_R   g2331( .A1 (x1), .A2 (n773), .B (n2338), .Y (y897) );
  AND3x1_ASAP7_75t_R   g2332( .A (n12), .B (x1), .C (x2), .Y (n2340) );
  INVx1_ASAP7_75t_R    g2333( .A (n2340), .Y (n2341) );
  AO32x1_ASAP7_75t_R   g2334( .A1 (n497), .A2 (n2341), .A3 (n746), .B1 (n15), .B2 (n1245), .Y (y898) );
  AO21x1_ASAP7_75t_R   g2335( .A1 (n436), .A2 (n466), .B (x5), .Y (n2343) );
  OA21x2_ASAP7_75t_R   g2336( .A1 (n537), .A2 (n463), .B (n2343), .Y (y899) );
  AND2x2_ASAP7_75t_R   g2337( .A (n1300), .B (n1646), .Y (n2345) );
  AO21x1_ASAP7_75t_R   g2338( .A1 (n1635), .A2 (y1356), .B (n2345), .Y (y900) );
  INVx1_ASAP7_75t_R    g2339( .A (n763), .Y (n2347) );
  AO21x1_ASAP7_75t_R   g2340( .A1 (n762), .A2 (n67), .B (n2347), .Y (y901) );
  AND2x2_ASAP7_75t_R   g2341( .A (n872), .B (n866), .Y (y902) );
  AND3x1_ASAP7_75t_R   g2342( .A (n2322), .B (n1562), .C (n1265), .Y (y903) );
  NAND2x1_ASAP7_75t_R  g2343( .A (x5), .B (n1257), .Y (n2351) );
  AO21x1_ASAP7_75t_R   g2344( .A1 (n2351), .A2 (n244), .B (n826), .Y (y904) );
  AO21x1_ASAP7_75t_R   g2345( .A1 (n1614), .A2 (x0), .B (n2122), .Y (y905) );
  AO32x1_ASAP7_75t_R   g2346( .A1 (n244), .A2 (n2351), .A3 (n827), .B1 (n15), .B2 (n1245), .Y (y906) );
  AO21x1_ASAP7_75t_R   g2347( .A1 (n765), .A2 (x1), .B (n1245), .Y (n2355) );
  INVx1_ASAP7_75t_R    g2348( .A (n2199), .Y (n2356) );
  AO21x1_ASAP7_75t_R   g2349( .A1 (n15), .A2 (n2355), .B (n2356), .Y (y907) );
  AO21x1_ASAP7_75t_R   g2350( .A1 (n64), .A2 (n63), .B (n12), .Y (n2358) );
  NOR2x1_ASAP7_75t_R   g2351( .A (y2079), .B (n2358), .Y (n2359) );
  INVx1_ASAP7_75t_R    g2352( .A (n2359), .Y (n2360) );
  AND2x2_ASAP7_75t_R   g2353( .A (n2360), .B (n1639), .Y (y908) );
  NAND2x1_ASAP7_75t_R  g2354( .A (n12), .B (n1529), .Y (n2362) );
  NOR2x1_ASAP7_75t_R   g2355( .A (x2), .B (n1092), .Y (n2363) );
  AO21x1_ASAP7_75t_R   g2356( .A1 (n497), .A2 (n2362), .B (n2363), .Y (n2364) );
  INVx1_ASAP7_75t_R    g2357( .A (n1529), .Y (n2365) );
  NAND2x1_ASAP7_75t_R  g2358( .A (n2365), .B (y772), .Y (n2366) );
  AND2x2_ASAP7_75t_R   g2359( .A (n2364), .B (n2366), .Y (y909) );
  OA211x2_ASAP7_75t_R  g2360( .A1 (n2365), .A2 (y772), .B (n2366), .C (y9), .Y (y910) );
  AND3x1_ASAP7_75t_R   g2361( .A (n219), .B (n90), .C (n15), .Y (n2369) );
  INVx1_ASAP7_75t_R    g2362( .A (n2369), .Y (n2370) );
  AND2x2_ASAP7_75t_R   g2363( .A (n2370), .B (n2182), .Y (y911) );
  AND3x1_ASAP7_75t_R   g2364( .A (n2322), .B (n2133), .C (n244), .Y (y912) );
  OA21x2_ASAP7_75t_R   g2365( .A1 (y772), .A2 (n1636), .B (n2133), .Y (y913) );
  AO21x1_ASAP7_75t_R   g2366( .A1 (n12), .A2 (n17), .B (y39), .Y (y914) );
  OR3x1_ASAP7_75t_R    g2367( .A (n848), .B (n495), .C (n61), .Y (y915) );
  AO33x2_ASAP7_75t_R   g2368( .A1 (x1), .A2 (x5), .A3 (n241), .B1 (n750), .B2 (n1624), .B3 (x0), .Y (y916) );
  AND2x2_ASAP7_75t_R   g2369( .A (n1912), .B (n2117), .Y (y917) );
  AND3x1_ASAP7_75t_R   g2370( .A (n90), .B (n219), .C (n2172), .Y (y1751) );
  AO21x1_ASAP7_75t_R   g2371( .A1 (n221), .A2 (n15), .B (y1751), .Y (y918) );
  AO32x1_ASAP7_75t_R   g2372( .A1 (n15), .A2 (n2162), .A3 (y9), .B1 (x2), .B2 (y873), .Y (y919) );
  AO21x1_ASAP7_75t_R   g2373( .A1 (n2210), .A2 (n16), .B (n1537), .Y (n2381) );
  XOR2x2_ASAP7_75t_R   g2374( .A (n2381), .B (x0), .Y (y920) );
  AO21x1_ASAP7_75t_R   g2375( .A1 (n174), .A2 (x5), .B (y435), .Y (n2383) );
  OA21x2_ASAP7_75t_R   g2376( .A1 (n2315), .A2 (n969), .B (n2383), .Y (y921) );
  AO21x1_ASAP7_75t_R   g2377( .A1 (x1), .A2 (n58), .B (n1762), .Y (y922) );
  AO32x1_ASAP7_75t_R   g2378( .A1 (n746), .A2 (x1), .A3 (n244), .B1 (n207), .B2 (y3852), .Y (y923) );
  AO21x1_ASAP7_75t_R   g2379( .A1 (n16), .A2 (n15), .B (n17), .Y (n2387) );
  AO21x1_ASAP7_75t_R   g2380( .A1 (n2387), .A2 (n1613), .B (y69), .Y (y924) );
  AO21x1_ASAP7_75t_R   g2381( .A1 (n232), .A2 (x2), .B (n1669), .Y (y925) );
  AND2x2_ASAP7_75t_R   g2382( .A (n1201), .B (n219), .Y (y926) );
  AO21x1_ASAP7_75t_R   g2383( .A1 (n16), .A2 (x2), .B (n544), .Y (n2391) );
  AO21x1_ASAP7_75t_R   g2384( .A1 (n2391), .A2 (n752), .B (n2329), .Y (y927) );
  NOR2x1_ASAP7_75t_R   g2385( .A (y2079), .B (n1490), .Y (n2393) );
  INVx1_ASAP7_75t_R    g2386( .A (n2393), .Y (n2394) );
  AND2x2_ASAP7_75t_R   g2387( .A (n2394), .B (n2282), .Y (y928) );
  OA21x2_ASAP7_75t_R   g2388( .A1 (n2038), .A2 (n969), .B (n2117), .Y (y929) );
  AND3x1_ASAP7_75t_R   g2389( .A (n12), .B (n15), .C (x5), .Y (n2397) );
  AO21x1_ASAP7_75t_R   g2390( .A1 (n97), .A2 (x0), .B (n2397), .Y (n2398) );
  AO21x1_ASAP7_75t_R   g2391( .A1 (n2398), .A2 (x1), .B (n732), .Y (y930) );
  OR3x1_ASAP7_75t_R    g2392( .A (y863), .B (y2079), .C (n22), .Y (y2250) );
  AND2x2_ASAP7_75t_R   g2393( .A (y2250), .B (n947), .Y (y931) );
  AND3x1_ASAP7_75t_R   g2394( .A (n1912), .B (n1639), .C (n64), .Y (y932) );
  AND2x2_ASAP7_75t_R   g2395( .A (y535), .B (n64), .Y (y933) );
  OR3x1_ASAP7_75t_R    g2396( .A (n43), .B (y2079), .C (x2), .Y (n2404) );
  INVx1_ASAP7_75t_R    g2397( .A (n2404), .Y (n2405) );
  OA21x2_ASAP7_75t_R   g2398( .A1 (n2405), .A2 (n143), .B (n1912), .Y (y934) );
  AO21x1_ASAP7_75t_R   g2399( .A1 (x1), .A2 (x0), .B (n15), .Y (n2407) );
  AND3x1_ASAP7_75t_R   g2400( .A (y6), .B (n1232), .C (n2407), .Y (y935) );
  AND3x1_ASAP7_75t_R   g2401( .A (n2116), .B (n2117), .C (y9), .Y (y936) );
  AND3x1_ASAP7_75t_R   g2402( .A (y855), .B (n228), .C (n17), .Y (n2410) );
  AO21x1_ASAP7_75t_R   g2403( .A1 (y855), .A2 (n228), .B (n17), .Y (n2411) );
  INVx1_ASAP7_75t_R    g2404( .A (n2411), .Y (n2412) );
  NOR2x1_ASAP7_75t_R   g2405( .A (n2410), .B (n2412), .Y (y937) );
  OR3x1_ASAP7_75t_R    g2406( .A (n211), .B (n16), .C (n12), .Y (n2414) );
  AO21x1_ASAP7_75t_R   g2407( .A1 (n15), .A2 (x0), .B (n17), .Y (n2415) );
  AO21x1_ASAP7_75t_R   g2408( .A1 (n244), .A2 (x1), .B (n2415), .Y (n2416) );
  AND2x2_ASAP7_75t_R   g2409( .A (n2414), .B (n2416), .Y (y938) );
  INVx1_ASAP7_75t_R    g2410( .A (n216), .Y (n2418) );
  AND3x1_ASAP7_75t_R   g2411( .A (n243), .B (x2), .C (x0), .Y (n2419) );
  AO21x1_ASAP7_75t_R   g2412( .A1 (n2418), .A2 (n175), .B (n2419), .Y (y940) );
  INVx1_ASAP7_75t_R    g2413( .A (n863), .Y (n2421) );
  OA21x2_ASAP7_75t_R   g2414( .A1 (n2421), .A2 (n1254), .B (n2416), .Y (y941) );
  AND3x1_ASAP7_75t_R   g2415( .A (n12), .B (x2), .C (x3), .Y (n2423) );
  INVx1_ASAP7_75t_R    g2416( .A (n2423), .Y (n2424) );
  AO32x1_ASAP7_75t_R   g2417( .A1 (n2424), .A2 (n2261), .A3 (n210), .B1 (n1838), .B2 (n1545), .Y (y942) );
  AND3x1_ASAP7_75t_R   g2418( .A (n2263), .B (n2271), .C (n228), .Y (y943) );
  INVx1_ASAP7_75t_R    g2419( .A (n1698), .Y (n2427) );
  AO32x1_ASAP7_75t_R   g2420( .A1 (n267), .A2 (n1698), .A3 (n1699), .B1 (n2427), .B2 (n16), .Y (y944) );
  AND3x1_ASAP7_75t_R   g2421( .A (n2273), .B (n2274), .C (n228), .Y (y945) );
  AO21x1_ASAP7_75t_R   g2422( .A1 (n482), .A2 (y195), .B (n306), .Y (y946) );
  AND3x1_ASAP7_75t_R   g2423( .A (n469), .B (n1720), .C (y9), .Y (y947) );
  AO21x1_ASAP7_75t_R   g2424( .A1 (n16), .A2 (n12), .B (n211), .Y (n2432) );
  AO21x1_ASAP7_75t_R   g2425( .A1 (n15), .A2 (n17), .B (y863), .Y (n2433) );
  AND2x2_ASAP7_75t_R   g2426( .A (n2432), .B (n2433), .Y (n2434) );
  AO21x1_ASAP7_75t_R   g2427( .A1 (n218), .A2 (n221), .B (n2434), .Y (y948) );
  OR3x1_ASAP7_75t_R    g2428( .A (n76), .B (n16), .C (n12), .Y (n2436) );
  AO21x1_ASAP7_75t_R   g2429( .A1 (y9), .A2 (n77), .B (n143), .Y (n2437) );
  AND3x1_ASAP7_75t_R   g2430( .A (n2436), .B (n2437), .C (n1572), .Y (y949) );
  AO21x1_ASAP7_75t_R   g2431( .A1 (x0), .A2 (n1510), .B (n54), .Y (y950) );
  INVx1_ASAP7_75t_R    g2432( .A (n1528), .Y (n2440) );
  AND3x1_ASAP7_75t_R   g2433( .A (x0), .B (x2), .C (x1), .Y (n2441) );
  OR3x1_ASAP7_75t_R    g2434( .A (n2440), .B (n53), .C (n2441), .Y (y951) );
  INVx1_ASAP7_75t_R    g2435( .A (n2391), .Y (n2443) );
  AO21x1_ASAP7_75t_R   g2436( .A1 (n497), .A2 (n276), .B (n2443), .Y (y952) );
  INVx1_ASAP7_75t_R    g2437( .A (n1106), .Y (n2445) );
  OR3x1_ASAP7_75t_R    g2438( .A (n2160), .B (n2445), .C (n1644), .Y (y953) );
  AO21x1_ASAP7_75t_R   g2439( .A1 (n352), .A2 (n128), .B (n495), .Y (n2447) );
  AO21x1_ASAP7_75t_R   g2440( .A1 (n276), .A2 (n497), .B (n2447), .Y (y954) );
  AO21x1_ASAP7_75t_R   g2441( .A1 (y2079), .A2 (x1), .B (n1644), .Y (n2449) );
  AO21x1_ASAP7_75t_R   g2442( .A1 (n276), .A2 (n497), .B (n2449), .Y (y955) );
  OA21x2_ASAP7_75t_R   g2443( .A1 (n1646), .A2 (y873), .B (n2116), .Y (y956) );
  AO21x1_ASAP7_75t_R   g2444( .A1 (y2079), .A2 (x0), .B (n128), .Y (n2452) );
  AO21x1_ASAP7_75t_R   g2445( .A1 (n989), .A2 (x2), .B (n2452), .Y (y957) );
  NAND2x1_ASAP7_75t_R  g2446( .A (n856), .B (n219), .Y (n2454) );
  INVx1_ASAP7_75t_R    g2447( .A (n1403), .Y (n2455) );
  AO21x1_ASAP7_75t_R   g2448( .A1 (x0), .A2 (x1), .B (n2455), .Y (n2456) );
  AND2x2_ASAP7_75t_R   g2449( .A (n2454), .B (n2456), .Y (y958) );
  INVx1_ASAP7_75t_R    g2450( .A (n1954), .Y (n2458) );
  OA33x2_ASAP7_75t_R   g2451( .A1 (n143), .A2 (n2458), .A3 (n15), .B1 (x2), .B2 (n481), .B3 (n1545), .Y (y959) );
  OR3x1_ASAP7_75t_R    g2452( .A (n2147), .B (y2196), .C (n1644), .Y (y960) );
  AO21x1_ASAP7_75t_R   g2453( .A1 (n556), .A2 (n228), .B (n1180), .Y (y961) );
  AND3x1_ASAP7_75t_R   g2454( .A (y2079), .B (x2), .C (x0), .Y (n2462) );
  INVx1_ASAP7_75t_R    g2455( .A (n1502), .Y (n2463) );
  OA33x2_ASAP7_75t_R   g2456( .A1 (n2462), .A2 (n989), .A3 (n2463), .B1 (n16), .B2 (x2), .B3 (y2196), .Y (y962) );
  AO21x1_ASAP7_75t_R   g2457( .A1 (n63), .A2 (n244), .B (y2079), .Y (n2465) );
  AND3x1_ASAP7_75t_R   g2458( .A (n16), .B (x2), .C (x0), .Y (n2466) );
  INVx1_ASAP7_75t_R    g2459( .A (n2466), .Y (n2467) );
  AND2x2_ASAP7_75t_R   g2460( .A (n2465), .B (n2467), .Y (y963) );
  AND3x1_ASAP7_75t_R   g2461( .A (n2116), .B (n2117), .C (n255), .Y (y964) );
  AO21x1_ASAP7_75t_R   g2462( .A1 (x0), .A2 (x2), .B (y2079), .Y (n2470) );
  NOR2x1_ASAP7_75t_R   g2463( .A (x1), .B (n2136), .Y (n2471) );
  AO21x1_ASAP7_75t_R   g2464( .A1 (n2470), .A2 (n747), .B (n2471), .Y (y965) );
  OR3x1_ASAP7_75t_R    g2465( .A (n2160), .B (n363), .C (n1644), .Y (y966) );
  AND2x2_ASAP7_75t_R   g2466( .A (n97), .B (n244), .Y (n2474) );
  INVx1_ASAP7_75t_R    g2467( .A (n2474), .Y (n2475) );
  OA21x2_ASAP7_75t_R   g2468( .A1 (n2475), .A2 (x1), .B (n2465), .Y (y967) );
  OR3x1_ASAP7_75t_R    g2469( .A (n2160), .B (n701), .C (n128), .Y (y968) );
  AO21x1_ASAP7_75t_R   g2470( .A1 (n12), .A2 (y2079), .B (n544), .Y (n2478) );
  INVx1_ASAP7_75t_R    g2471( .A (n2478), .Y (n2479) );
  AO32x1_ASAP7_75t_R   g2472( .A1 (y3852), .A2 (n90), .A3 (x2), .B1 (n2479), .B2 (n15), .Y (y969) );
  AO21x1_ASAP7_75t_R   g2473( .A1 (y2079), .A2 (x2), .B (n128), .Y (n2481) );
  AO21x1_ASAP7_75t_R   g2474( .A1 (n352), .A2 (n2481), .B (n2160), .Y (y970) );
  AND3x1_ASAP7_75t_R   g2475( .A (n90), .B (n219), .C (y2079), .Y (y2219) );
  OA33x2_ASAP7_75t_R   g2476( .A1 (n15), .A2 (n495), .A3 (y772), .B1 (x2), .B2 (n1259), .B3 (y2219), .Y (y971) );
  OR3x1_ASAP7_75t_R    g2477( .A (n2441), .B (n363), .C (n51), .Y (y972) );
  AO21x1_ASAP7_75t_R   g2478( .A1 (n1910), .A2 (n63), .B (n363), .Y (y973) );
  AND2x2_ASAP7_75t_R   g2479( .A (y972), .B (n93), .Y (y974) );
  AO21x1_ASAP7_75t_R   g2480( .A1 (n2470), .A2 (x1), .B (n2471), .Y (y975) );
  NAND2x1_ASAP7_75t_R  g2481( .A (n16), .B (n1502), .Y (n2489) );
  OR3x1_ASAP7_75t_R    g2482( .A (n276), .B (y2079), .C (n16), .Y (n2490) );
  AND2x2_ASAP7_75t_R   g2483( .A (n2489), .B (n2490), .Y (y976) );
  AO21x1_ASAP7_75t_R   g2484( .A1 (n16), .A2 (n15), .B (n1503), .Y (y977) );
  AO21x1_ASAP7_75t_R   g2485( .A1 (n12), .A2 (y2079), .B (n276), .Y (n2493) );
  OA21x2_ASAP7_75t_R   g2486( .A1 (n2493), .A2 (n16), .B (n64), .Y (y978) );
  AO21x1_ASAP7_75t_R   g2487( .A1 (n352), .A2 (n128), .B (n2147), .Y (y979) );
  AND3x1_ASAP7_75t_R   g2488( .A (n497), .B (n219), .C (x2), .Y (n2496) );
  AO21x1_ASAP7_75t_R   g2489( .A1 (n15), .A2 (n776), .B (n2496), .Y (y980) );
  NAND2x1_ASAP7_75t_R  g2490( .A (n994), .B (n312), .Y (n2498) );
  AO21x1_ASAP7_75t_R   g2491( .A1 (n2498), .A2 (n15), .B (n2496), .Y (y981) );
  AO32x1_ASAP7_75t_R   g2492( .A1 (n12), .A2 (n63), .A3 (n497), .B1 (x5), .B2 (n2326), .Y (n2500) );
  INVx1_ASAP7_75t_R    g2493( .A (n2500), .Y (y982) );
  AO21x1_ASAP7_75t_R   g2494( .A1 (n2208), .A2 (n758), .B (n2169), .Y (y983) );
  AO21x1_ASAP7_75t_R   g2495( .A1 (n15), .A2 (x5), .B (x1), .Y (n2503) );
  INVx1_ASAP7_75t_R    g2496( .A (n2503), .Y (n2504) );
  AOI22x1_ASAP7_75t_R  g2497( .A1 (n2504), .A2 (n1387), .B1 (n2475), .B2 (x1), .Y (y984) );
  AO21x1_ASAP7_75t_R   g2498( .A1 (n16), .A2 (n2208), .B (n2160), .Y (y985) );
  INVx1_ASAP7_75t_R    g2499( .A (n2095), .Y (n2507) );
  INVx1_ASAP7_75t_R    g2500( .A (n1542), .Y (n2508) );
  OR3x1_ASAP7_75t_R    g2501( .A (n363), .B (n15), .C (x1), .Y (n2509) );
  OA21x2_ASAP7_75t_R   g2502( .A1 (n2507), .A2 (n2508), .B (n2509), .Y (y986) );
  AO21x1_ASAP7_75t_R   g2503( .A1 (n12), .A2 (x1), .B (x2), .Y (n2511) );
  OA22x2_ASAP7_75t_R   g2504( .A1 (n2511), .A2 (n1245), .B1 (y1356), .B2 (n15), .Y (y987) );
  AO21x1_ASAP7_75t_R   g2505( .A1 (y2079), .A2 (x0), .B (n756), .Y (n2513) );
  INVx1_ASAP7_75t_R    g2506( .A (n2513), .Y (n2514) );
  OA22x2_ASAP7_75t_R   g2507( .A1 (n16), .A2 (n2513), .B1 (n143), .B2 (n2514), .Y (y988) );
  NAND2x1_ASAP7_75t_R  g2508( .A (n1510), .B (n65), .Y (n2516) );
  OA21x2_ASAP7_75t_R   g2509( .A1 (n694), .A2 (n1525), .B (n2516), .Y (y989) );
  NAND2x1_ASAP7_75t_R  g2510( .A (n750), .B (n64), .Y (n2518) );
  AOI21x1_ASAP7_75t_R  g2511( .A1 (n583), .A2 (n2518), .B (n2340), .Y (y990) );
  NOR2x1_ASAP7_75t_R   g2512( .A (n43), .B (n1696), .Y (y991) );
  AND2x2_ASAP7_75t_R   g2513( .A (n1640), .B (n2117), .Y (y992) );
  AO21x1_ASAP7_75t_R   g2514( .A1 (n15), .A2 (y9), .B (n1910), .Y (n2522) );
  AND2x2_ASAP7_75t_R   g2515( .A (n2522), .B (n1640), .Y (y993) );
  AO21x1_ASAP7_75t_R   g2516( .A1 (x5), .A2 (n15), .B (n90), .Y (n2524) );
  AND3x1_ASAP7_75t_R   g2517( .A (n2524), .B (n1640), .C (n244), .Y (y994) );
  AND2x2_ASAP7_75t_R   g2518( .A (n895), .B (x0), .Y (y995) );
  AND3x1_ASAP7_75t_R   g2519( .A (n97), .B (n244), .C (x1), .Y (n2527) );
  AO21x1_ASAP7_75t_R   g2520( .A1 (n16), .A2 (n1646), .B (n2527), .Y (y996) );
  AO21x1_ASAP7_75t_R   g2521( .A1 (n1643), .A2 (x0), .B (n128), .Y (y997) );
  AO21x1_ASAP7_75t_R   g2522( .A1 (n352), .A2 (n128), .B (n2160), .Y (y998) );
  AO21x1_ASAP7_75t_R   g2523( .A1 (n1643), .A2 (x0), .B (n1644), .Y (y999) );
  OR3x1_ASAP7_75t_R    g2524( .A (n363), .B (n16), .C (x2), .Y (n2532) );
  AND2x2_ASAP7_75t_R   g2525( .A (n2532), .B (n2117), .Y (y1000) );
  AND2x2_ASAP7_75t_R   g2526( .A (n776), .B (n352), .Y (n2534) );
  OA21x2_ASAP7_75t_R   g2527( .A1 (n2534), .A2 (x2), .B (n2117), .Y (y1001) );
  AND3x1_ASAP7_75t_R   g2528( .A (n64), .B (n63), .C (n1480), .Y (y1002) );
  AO21x1_ASAP7_75t_R   g2529( .A1 (n125), .A2 (n51), .B (n2441), .Y (y1003) );
  AO21x1_ASAP7_75t_R   g2530( .A1 (n15), .A2 (x3), .B (n143), .Y (n2538) );
  AND2x2_ASAP7_75t_R   g2531( .A (n2538), .B (n63), .Y (y1004) );
  INVx1_ASAP7_75t_R    g2532( .A (n913), .Y (n2540) );
  AO21x1_ASAP7_75t_R   g2533( .A1 (y2079), .A2 (n63), .B (n2540), .Y (y1005) );
  INVx1_ASAP7_75t_R    g2534( .A (n1029), .Y (n2542) );
  AND2x2_ASAP7_75t_R   g2535( .A (n496), .B (n2542), .Y (y1006) );
  AND3x1_ASAP7_75t_R   g2536( .A (n145), .B (x1), .C (x2), .Y (n2544) );
  AO21x1_ASAP7_75t_R   g2537( .A1 (n15), .A2 (n16), .B (n139), .Y (n2545) );
  INVx1_ASAP7_75t_R    g2538( .A (n878), .Y (n2546) );
  OR3x1_ASAP7_75t_R    g2539( .A (n2544), .B (n2545), .C (n2546), .Y (y1007) );
  NAND2x1_ASAP7_75t_R  g2540( .A (n51), .B (n125), .Y (n2548) );
  INVx1_ASAP7_75t_R    g2541( .A (n2441), .Y (n2549) );
  AO32x1_ASAP7_75t_R   g2542( .A1 (n2548), .A2 (n2549), .A3 (n17), .B1 (x3), .B2 (y1003), .Y (y1008) );
  NAND2x1_ASAP7_75t_R  g2543( .A (n2158), .B (n64), .Y (n2551) );
  AO21x1_ASAP7_75t_R   g2544( .A1 (n64), .A2 (n2158), .B (n17), .Y (n2552) );
  OA21x2_ASAP7_75t_R   g2545( .A1 (n2551), .A2 (x3), .B (n2552), .Y (y3143) );
  AO21x1_ASAP7_75t_R   g2546( .A1 (n12), .A2 (n17), .B (y3143), .Y (y1009) );
  AO21x1_ASAP7_75t_R   g2547( .A1 (x0), .A2 (x2), .B (x3), .Y (n2555) );
  INVx1_ASAP7_75t_R    g2548( .A (n2555), .Y (n2556) );
  AO21x1_ASAP7_75t_R   g2549( .A1 (x2), .A2 (n145), .B (n2556), .Y (n2557) );
  AO22x1_ASAP7_75t_R   g2550( .A1 (n16), .A2 (n863), .B1 (x1), .B2 (n2557), .Y (y1010) );
  NAND2x1_ASAP7_75t_R  g2551( .A (n2117), .B (n63), .Y (n2559) );
  AO21x1_ASAP7_75t_R   g2552( .A1 (n12), .A2 (n16), .B (x3), .Y (n2560) );
  XOR2x2_ASAP7_75t_R   g2553( .A (n2559), .B (n2560), .Y (y1011) );
  AO21x1_ASAP7_75t_R   g2554( .A1 (n17), .A2 (y25), .B (n2441), .Y (n2562) );
  NAND2x1_ASAP7_75t_R  g2555( .A (x0), .B (n235), .Y (n2563) );
  OA21x2_ASAP7_75t_R   g2556( .A1 (n51), .A2 (n2562), .B (n2563), .Y (y1012) );
  AND3x1_ASAP7_75t_R   g2557( .A (x0), .B (x1), .C (x3), .Y (n2565) );
  INVx1_ASAP7_75t_R    g2558( .A (n2565), .Y (n2566) );
  AO21x1_ASAP7_75t_R   g2559( .A1 (n219), .A2 (n90), .B (x3), .Y (n2567) );
  AO21x1_ASAP7_75t_R   g2560( .A1 (n125), .A2 (x1), .B (n122), .Y (n2568) );
  AO32x1_ASAP7_75t_R   g2561( .A1 (x2), .A2 (n2566), .A3 (n2567), .B1 (n15), .B2 (n2568), .Y (n2569) );
  INVx1_ASAP7_75t_R    g2562( .A (n2569), .Y (y1013) );
  NAND2x1_ASAP7_75t_R  g2563( .A (n328), .B (n382), .Y (n2571) );
  AND3x1_ASAP7_75t_R   g2564( .A (n12), .B (x3), .C (x5), .Y (n2572) );
  NAND2x1_ASAP7_75t_R  g2565( .A (x4), .B (n2572), .Y (n2573) );
  OA21x2_ASAP7_75t_R   g2566( .A1 (n2571), .A2 (n481), .B (n2573), .Y (y1014) );
  AO21x1_ASAP7_75t_R   g2567( .A1 (n17), .A2 (x1), .B (n15), .Y (n2575) );
  AND3x1_ASAP7_75t_R   g2568( .A (n17), .B (x1), .C (x0), .Y (n2576) );
  INVx1_ASAP7_75t_R    g2569( .A (n2576), .Y (n2577) );
  AO21x1_ASAP7_75t_R   g2570( .A1 (n16), .A2 (x3), .B (n2576), .Y (n2578) );
  AO32x1_ASAP7_75t_R   g2571( .A1 (n1296), .A2 (n2577), .A3 (x2), .B1 (n15), .B2 (n2578), .Y (n2579) );
  OA21x2_ASAP7_75t_R   g2572( .A1 (x0), .A2 (n2575), .B (n2579), .Y (y1015) );
  AND3x1_ASAP7_75t_R   g2573( .A (n145), .B (x2), .C (x1), .Y (n2581) );
  OR3x1_ASAP7_75t_R    g2574( .A (n2581), .B (n2556), .C (n128), .Y (y1016) );
  INVx1_ASAP7_75t_R    g2575( .A (n1301), .Y (n2583) );
  AO32x1_ASAP7_75t_R   g2576( .A1 (n84), .A2 (n2583), .A3 (n125), .B1 (n15), .B2 (n611), .Y (y1017) );
  AO21x1_ASAP7_75t_R   g2577( .A1 (n12), .A2 (n17), .B (n243), .Y (n2585) );
  AOI22x1_ASAP7_75t_R  g2578( .A1 (n15), .A2 (n2585), .B1 (n203), .B2 (n2566), .Y (y1018) );
  AO21x1_ASAP7_75t_R   g2579( .A1 (n17), .A2 (x2), .B (n128), .Y (n2587) );
  NOR2x1_ASAP7_75t_R   g2580( .A (n105), .B (n133), .Y (n2588) );
  AO21x1_ASAP7_75t_R   g2581( .A1 (n125), .A2 (n2587), .B (n2588), .Y (y1019) );
  AND3x1_ASAP7_75t_R   g2582( .A (x0), .B (x2), .C (x3), .Y (n2590) );
  AO21x1_ASAP7_75t_R   g2583( .A1 (x1), .A2 (n2590), .B (n2545), .Y (y1020) );
  AO21x1_ASAP7_75t_R   g2584( .A1 (n2542), .A2 (n299), .B (y2079), .Y (y1021) );
  AND2x2_ASAP7_75t_R   g2585( .A (n64), .B (n1635), .Y (n2593) );
  AO21x1_ASAP7_75t_R   g2586( .A1 (n2549), .A2 (n52), .B (n17), .Y (n2594) );
  OAI21x1_ASAP7_75t_R  g2587( .A1 (x3), .A2 (n2593), .B (n2594), .Y (y1022) );
  NAND2x1_ASAP7_75t_R  g2588( .A (n43), .B (n28), .Y (n2596) );
  INVx1_ASAP7_75t_R    g2589( .A (n2596), .Y (n2597) );
  AO21x1_ASAP7_75t_R   g2590( .A1 (n2597), .A2 (n447), .B (y1775), .Y (y1023) );
  AO21x1_ASAP7_75t_R   g2591( .A1 (n1564), .A2 (n63), .B (y2079), .Y (y1024) );
  NOR2x1_ASAP7_75t_R   g2592( .A (x5), .B (n330), .Y (n2600) );
  AO21x1_ASAP7_75t_R   g2593( .A1 (n1791), .A2 (n652), .B (n2600), .Y (y1025) );
  NOR2x1_ASAP7_75t_R   g2594( .A (n1450), .B (n610), .Y (n2602) );
  AO21x1_ASAP7_75t_R   g2595( .A1 (y2079), .A2 (n827), .B (n2602), .Y (y1026) );
  AND2x2_ASAP7_75t_R   g2596( .A (y1024), .B (n93), .Y (y1027) );
  NAND2x1_ASAP7_75t_R  g2597( .A (x5), .B (n610), .Y (n2605) );
  AND2x2_ASAP7_75t_R   g2598( .A (n2605), .B (n2307), .Y (y1028) );
  AO21x1_ASAP7_75t_R   g2599( .A1 (x2), .A2 (x5), .B (n12), .Y (n2607) );
  NAND2x1_ASAP7_75t_R  g2600( .A (n16), .B (n2607), .Y (n2608) );
  AND2x2_ASAP7_75t_R   g2601( .A (n2608), .B (n2490), .Y (y1029) );
  AND2x2_ASAP7_75t_R   g2602( .A (n750), .B (x0), .Y (n2610) );
  OA21x2_ASAP7_75t_R   g2603( .A1 (n590), .A2 (n2610), .B (n2307), .Y (y1030) );
  OR3x1_ASAP7_75t_R    g2604( .A (n2397), .B (n16), .C (n276), .Y (n2612) );
  OA21x2_ASAP7_75t_R   g2605( .A1 (n363), .A2 (n851), .B (n2612), .Y (y1031) );
  AO21x1_ASAP7_75t_R   g2606( .A1 (y2079), .A2 (y1116), .B (y2259), .Y (y1032) );
  AO21x1_ASAP7_75t_R   g2607( .A1 (n1176), .A2 (x5), .B (n1004), .Y (y1033) );
  AND2x2_ASAP7_75t_R   g2608( .A (n2605), .B (n2467), .Y (y1034) );
  AND2x2_ASAP7_75t_R   g2609( .A (n2605), .B (n2524), .Y (y1035) );
  OA21x2_ASAP7_75t_R   g2610( .A1 (n2475), .A2 (x1), .B (n2605), .Y (y1036) );
  AO21x1_ASAP7_75t_R   g2611( .A1 (n1352), .A2 (n15), .B (n2466), .Y (n2619) );
  NOR2x1_ASAP7_75t_R   g2612( .A (n481), .B (n2619), .Y (y1037) );
  AND2x2_ASAP7_75t_R   g2613( .A (n740), .B (n90), .Y (n2621) );
  AOI21x1_ASAP7_75t_R  g2614( .A1 (n1542), .A2 (n2621), .B (n2466), .Y (y1038) );
  NAND2x1_ASAP7_75t_R  g2615( .A (n15), .B (n1352), .Y (n2623) );
  AND3x1_ASAP7_75t_R   g2616( .A (n2623), .B (n2524), .C (y3852), .Y (y1039) );
  AND3x1_ASAP7_75t_R   g2617( .A (n64), .B (n750), .C (x0), .Y (n2625) );
  AO21x1_ASAP7_75t_R   g2618( .A1 (n12), .A2 (y2079), .B (n2625), .Y (y1040) );
  NAND2x1_ASAP7_75t_R  g2619( .A (n93), .B (n155), .Y (y1762) );
  AOI21x1_ASAP7_75t_R  g2620( .A1 (n14), .A2 (y1762), .B (n481), .Y (y1041) );
  INVx1_ASAP7_75t_R    g2621( .A (n1033), .Y (n2629) );
  AO21x1_ASAP7_75t_R   g2622( .A1 (n211), .A2 (x1), .B (x0), .Y (n2630) );
  AND2x2_ASAP7_75t_R   g2623( .A (n2629), .B (n2630), .Y (y1042) );
  AND2x2_ASAP7_75t_R   g2624( .A (n2605), .B (n64), .Y (y1043) );
  AO21x1_ASAP7_75t_R   g2625( .A1 (n1480), .A2 (n747), .B (n45), .Y (y1044) );
  OR3x1_ASAP7_75t_R    g2626( .A (n495), .B (n2169), .C (n826), .Y (y1045) );
  AND2x2_ASAP7_75t_R   g2627( .A (y3134), .B (n684), .Y (y1046) );
  OA21x2_ASAP7_75t_R   g2628( .A1 (n1682), .A2 (n1689), .B (n1690), .Y (y1047) );
  AND2x2_ASAP7_75t_R   g2629( .A (n2489), .B (n2605), .Y (y1048) );
  AO21x1_ASAP7_75t_R   g2630( .A1 (n2287), .A2 (n15), .B (n2147), .Y (y1049) );
  NAND2x1_ASAP7_75t_R  g2631( .A (n128), .B (n352), .Y (n2639) );
  INVx1_ASAP7_75t_R    g2632( .A (n2639), .Y (n2640) );
  AO21x1_ASAP7_75t_R   g2633( .A1 (n1502), .A2 (x1), .B (n2640), .Y (n2641) );
  AND2x2_ASAP7_75t_R   g2634( .A (n2641), .B (y3852), .Y (y1050) );
  AO21x1_ASAP7_75t_R   g2635( .A1 (n97), .A2 (x1), .B (n1644), .Y (n2643) );
  AND2x2_ASAP7_75t_R   g2636( .A (n2643), .B (n707), .Y (y1051) );
  AO21x1_ASAP7_75t_R   g2637( .A1 (x0), .A2 (x4), .B (x3), .Y (n2645) );
  OA21x2_ASAP7_75t_R   g2638( .A1 (n481), .A2 (n2645), .B (n922), .Y (y1052) );
  INVx1_ASAP7_75t_R    g2639( .A (n746), .Y (n2647) );
  OA21x2_ASAP7_75t_R   g2640( .A1 (n2647), .A2 (n989), .B (n2116), .Y (y1053) );
  AND3x1_ASAP7_75t_R   g2641( .A (n63), .B (y3852), .C (n64), .Y (y1054) );
  AO21x1_ASAP7_75t_R   g2642( .A1 (x5), .A2 (n12), .B (n64), .Y (n2650) );
  OA21x2_ASAP7_75t_R   g2643( .A1 (n1545), .A2 (n2210), .B (n2650), .Y (y1055) );
  NAND2x1_ASAP7_75t_R  g2644( .A (n15), .B (n994), .Y (n2652) );
  AND3x1_ASAP7_75t_R   g2645( .A (n2652), .B (n64), .C (y3852), .Y (y1056) );
  AND3x1_ASAP7_75t_R   g2646( .A (n64), .B (y3852), .C (n750), .Y (y1057) );
  AO21x1_ASAP7_75t_R   g2647( .A1 (n352), .A2 (n128), .B (n1503), .Y (y1058) );
  AO21x1_ASAP7_75t_R   g2648( .A1 (n694), .A2 (n1675), .B (n1464), .Y (y1059) );
  AO21x1_ASAP7_75t_R   g2649( .A1 (n16), .A2 (y2079), .B (n12), .Y (n2657) );
  INVx1_ASAP7_75t_R    g2650( .A (n2657), .Y (n2658) );
  OA21x2_ASAP7_75t_R   g2651( .A1 (n1676), .A2 (n2658), .B (n1586), .Y (y1060) );
  AND2x2_ASAP7_75t_R   g2652( .A (n2182), .B (n2211), .Y (y1061) );
  AO21x1_ASAP7_75t_R   g2653( .A1 (n15), .A2 (x1), .B (x0), .Y (n2661) );
  AND2x2_ASAP7_75t_R   g2654( .A (n1614), .B (n2661), .Y (y1062) );
  OR3x1_ASAP7_75t_R    g2655( .A (n1210), .B (n589), .C (x2), .Y (n2663) );
  NAND2x1_ASAP7_75t_R  g2656( .A (n2199), .B (n2663), .Y (y1063) );
  AO21x1_ASAP7_75t_R   g2657( .A1 (y2079), .A2 (x1), .B (n1245), .Y (n2665) );
  AO21x1_ASAP7_75t_R   g2658( .A1 (n2665), .A2 (n15), .B (n2356), .Y (y1064) );
  OA21x2_ASAP7_75t_R   g2659( .A1 (n978), .A2 (n2182), .B (n1912), .Y (y1065) );
  INVx1_ASAP7_75t_R    g2660( .A (n2140), .Y (n2668) );
  AND2x2_ASAP7_75t_R   g2661( .A (n1510), .B (x0), .Y (y1199) );
  AO21x1_ASAP7_75t_R   g2662( .A1 (n16), .A2 (n2668), .B (y1199), .Y (y1066) );
  AND3x1_ASAP7_75t_R   g2663( .A (n497), .B (n1529), .C (x0), .Y (y1201) );
  AO21x1_ASAP7_75t_R   g2664( .A1 (n988), .A2 (n2463), .B (y1201), .Y (n2672) );
  AND2x2_ASAP7_75t_R   g2665( .A (n2672), .B (y3852), .Y (y1068) );
  AO21x1_ASAP7_75t_R   g2666( .A1 (n16), .A2 (x0), .B (n103), .Y (n2674) );
  AO21x1_ASAP7_75t_R   g2667( .A1 (n219), .A2 (n90), .B (n15), .Y (n2675) );
  OA21x2_ASAP7_75t_R   g2668( .A1 (y2079), .A2 (n2674), .B (n2675), .Y (y1070) );
  OA21x2_ASAP7_75t_R   g2669( .A1 (n1087), .A2 (y195), .B (n968), .Y (y1071) );
  AO21x1_ASAP7_75t_R   g2670( .A1 (n2475), .A2 (n2317), .B (n2527), .Y (y1072) );
  INVx1_ASAP7_75t_R    g2671( .A (n103), .Y (n2679) );
  AO21x1_ASAP7_75t_R   g2672( .A1 (n847), .A2 (n2679), .B (n2169), .Y (y1073) );
  OA21x2_ASAP7_75t_R   g2673( .A1 (n559), .A2 (n2315), .B (n2467), .Y (y1074) );
  AND2x2_ASAP7_75t_R   g2674( .A (n1863), .B (y109), .Y (y1075) );
  AND3x1_ASAP7_75t_R   g2675( .A (n2605), .B (n1424), .C (n2467), .Y (y1076) );
  AO21x1_ASAP7_75t_R   g2676( .A1 (n77), .A2 (n674), .B (n12), .Y (n2684) );
  NAND2x1_ASAP7_75t_R  g2677( .A (n167), .B (n2684), .Y (y1077) );
  OA21x2_ASAP7_75t_R   g2678( .A1 (n559), .A2 (n2315), .B (n2524), .Y (y1078) );
  AO21x1_ASAP7_75t_R   g2679( .A1 (n1564), .A2 (n63), .B (n854), .Y (y1079) );
  NAND2x1_ASAP7_75t_R  g2680( .A (n12), .B (n763), .Y (n2688) );
  OA21x2_ASAP7_75t_R   g2681( .A1 (n53), .A2 (n703), .B (n2688), .Y (y1080) );
  OA21x2_ASAP7_75t_R   g2682( .A1 (n241), .A2 (n1910), .B (n2211), .Y (y1082) );
  AO21x1_ASAP7_75t_R   g2683( .A1 (n22), .A2 (n316), .B (n538), .Y (y1083) );
  AO21x1_ASAP7_75t_R   g2684( .A1 (n481), .A2 (n527), .B (n957), .Y (y1085) );
  AND2x2_ASAP7_75t_R   g2685( .A (n2503), .B (x0), .Y (n2693) );
  AO21x1_ASAP7_75t_R   g2686( .A1 (n2693), .A2 (n1640), .B (n2047), .Y (y1086) );
  AO21x1_ASAP7_75t_R   g2687( .A1 (n527), .A2 (n12), .B (n1809), .Y (y1087) );
  AO22x1_ASAP7_75t_R   g2688( .A1 (x1), .A2 (n1047), .B1 (n16), .B2 (n510), .Y (y1088) );
  AND2x2_ASAP7_75t_R   g2689( .A (n2643), .B (x0), .Y (y1089) );
  AO21x1_ASAP7_75t_R   g2690( .A1 (y3852), .A2 (n1454), .B (n2169), .Y (y1090) );
  AO21x1_ASAP7_75t_R   g2691( .A1 (n495), .A2 (n15), .B (x0), .Y (n2699) );
  AND2x2_ASAP7_75t_R   g2692( .A (n2699), .B (n2358), .Y (y1091) );
  AO21x1_ASAP7_75t_R   g2693( .A1 (x5), .A2 (n16), .B (n746), .Y (n2701) );
  OA21x2_ASAP7_75t_R   g2694( .A1 (n2647), .A2 (n1416), .B (n2701), .Y (y1092) );
  OA211x2_ASAP7_75t_R  g2695( .A1 (n1545), .A2 (n2136), .B (n2117), .C (n743), .Y (y1093) );
  AND3x1_ASAP7_75t_R   g2696( .A (n63), .B (n64), .C (n1066), .Y (y1094) );
  AND3x1_ASAP7_75t_R   g2697( .A (n145), .B (n15), .C (n16), .Y (n2705) );
  AO21x1_ASAP7_75t_R   g2698( .A1 (n210), .A2 (n746), .B (n2705), .Y (n2706) );
  AND2x2_ASAP7_75t_R   g2699( .A (n2706), .B (n219), .Y (y1095) );
  AND3x1_ASAP7_75t_R   g2700( .A (n64), .B (n1546), .C (x0), .Y (y1096) );
  AO21x1_ASAP7_75t_R   g2701( .A1 (n510), .A2 (n512), .B (n143), .Y (y1097) );
  INVx1_ASAP7_75t_R    g2702( .A (n611), .Y (n2710) );
  OR3x1_ASAP7_75t_R    g2703( .A (n2710), .B (n15), .C (n122), .Y (n2711) );
  AO21x1_ASAP7_75t_R   g2704( .A1 (x0), .A2 (n17), .B (n63), .Y (n2712) );
  AND3x1_ASAP7_75t_R   g2705( .A (n2711), .B (n2712), .C (n84), .Y (y1098) );
  INVx1_ASAP7_75t_R    g2706( .A (n25), .Y (n2714) );
  INVx1_ASAP7_75t_R    g2707( .A (n23), .Y (n2715) );
  AO21x1_ASAP7_75t_R   g2708( .A1 (n2714), .A2 (n2715), .B (n143), .Y (n2716) );
  AO21x1_ASAP7_75t_R   g2709( .A1 (y9), .A2 (y3758), .B (n2716), .Y (y1099) );
  INVx1_ASAP7_75t_R    g2710( .A (n125), .Y (n2718) );
  AND3x1_ASAP7_75t_R   g2711( .A (n2718), .B (n63), .C (n64), .Y (n2719) );
  INVx1_ASAP7_75t_R    g2712( .A (n2719), .Y (n2720) );
  AO21x1_ASAP7_75t_R   g2713( .A1 (n2315), .A2 (n64), .B (n17), .Y (n2721) );
  AO21x1_ASAP7_75t_R   g2714( .A1 (n64), .A2 (n63), .B (x0), .Y (n2722) );
  AND3x1_ASAP7_75t_R   g2715( .A (n2720), .B (n2721), .C (n2722), .Y (y1100) );
  AND2x2_ASAP7_75t_R   g2716( .A (n948), .B (x5), .Y (n2724) );
  AO221x2_ASAP7_75t_R  g2717( .A1 (n529), .A2 (n228), .B1 (n947), .B2 (n2724), .C (y863), .Y (y1101) );
  AO21x1_ASAP7_75t_R   g2718( .A1 (n17), .A2 (x1), .B (x0), .Y (n2726) );
  AND2x2_ASAP7_75t_R   g2719( .A (n2579), .B (n2726), .Y (y1102) );
  NAND2x1_ASAP7_75t_R  g2720( .A (x3), .B (n610), .Y (n2728) );
  OR3x1_ASAP7_75t_R    g2721( .A (n243), .B (n15), .C (n12), .Y (n2729) );
  AND2x2_ASAP7_75t_R   g2722( .A (n2728), .B (n2729), .Y (y1103) );
  AO21x1_ASAP7_75t_R   g2723( .A1 (n16), .A2 (x2), .B (n17), .Y (n2731) );
  NOR2x1_ASAP7_75t_R   g2724( .A (n2731), .B (n610), .Y (n2732) );
  AO21x1_ASAP7_75t_R   g2725( .A1 (n17), .A2 (n610), .B (n2732), .Y (y1104) );
  INVx1_ASAP7_75t_R    g2726( .A (n1297), .Y (n2734) );
  OA211x2_ASAP7_75t_R  g2727( .A1 (n2734), .A2 (x2), .B (n84), .C (n2729), .Y (y1105) );
  NAND2x1_ASAP7_75t_R  g2728( .A (n15), .B (n2710), .Y (n2736) );
  AND3x1_ASAP7_75t_R   g2729( .A (n2736), .B (n2729), .C (n84), .Y (y1106) );
  AO21x1_ASAP7_75t_R   g2730( .A1 (n15), .A2 (x3), .B (n12), .Y (n2738) );
  AND2x2_ASAP7_75t_R   g2731( .A (n137), .B (n90), .Y (n2739) );
  INVx1_ASAP7_75t_R    g2732( .A (n2729), .Y (n2740) );
  AOI21x1_ASAP7_75t_R  g2733( .A1 (n2738), .A2 (n2739), .B (n2740), .Y (y1107) );
  AO21x1_ASAP7_75t_R   g2734( .A1 (n17), .A2 (x2), .B (n16), .Y (n2742) );
  NAND2x1_ASAP7_75t_R  g2735( .A (n2738), .B (n2742), .Y (n2743) );
  INVx1_ASAP7_75t_R    g2736( .A (n2588), .Y (n2744) );
  AOI21x1_ASAP7_75t_R  g2737( .A1 (n2743), .A2 (n2744), .B (n1032), .Y (y1108) );
  INVx1_ASAP7_75t_R    g2738( .A (n2738), .Y (n2746) );
  OA33x2_ASAP7_75t_R   g2739( .A1 (n163), .A2 (n1545), .A3 (n2746), .B1 (n12), .B2 (n2739), .B3 (n164), .Y (y1109) );
  AO21x1_ASAP7_75t_R   g2740( .A1 (x2), .A2 (x3), .B (n16), .Y (n2748) );
  INVx1_ASAP7_75t_R    g2741( .A (n2748), .Y (n2749) );
  OR3x1_ASAP7_75t_R    g2742( .A (n1262), .B (n12), .C (n2749), .Y (n2750) );
  NAND2x1_ASAP7_75t_R  g2743( .A (n189), .B (n2750), .Y (y1111) );
  NAND2x1_ASAP7_75t_R  g2744( .A (n2748), .B (n64), .Y (n2752) );
  INVx1_ASAP7_75t_R    g2745( .A (n2752), .Y (n2753) );
  NAND2x1_ASAP7_75t_R  g2746( .A (n12), .B (n148), .Y (n2754) );
  OA21x2_ASAP7_75t_R   g2747( .A1 (n2753), .A2 (n12), .B (n2754), .Y (y1112) );
  AO21x1_ASAP7_75t_R   g2748( .A1 (n15), .A2 (x1), .B (n17), .Y (n2756) );
  INVx1_ASAP7_75t_R    g2749( .A (n2756), .Y (n2757) );
  AO21x1_ASAP7_75t_R   g2750( .A1 (n2757), .A2 (n1564), .B (n139), .Y (y1113) );
  INVx1_ASAP7_75t_R    g2751( .A (n176), .Y (y1114) );
  NAND2x1_ASAP7_75t_R  g2752( .A (n15), .B (n611), .Y (n2760) );
  NAND2x1_ASAP7_75t_R  g2753( .A (x1), .B (n2421), .Y (n2761) );
  AOI21x1_ASAP7_75t_R  g2754( .A1 (n2760), .A2 (n2761), .B (n1032), .Y (y1115) );
  AND3x1_ASAP7_75t_R   g2755( .A (n12), .B (n17), .C (x1), .Y (n2763) );
  AO32x1_ASAP7_75t_R   g2756( .A1 (n253), .A2 (n1554), .A3 (x0), .B1 (x2), .B2 (n2763), .Y (y1117) );
  AND3x1_ASAP7_75t_R   g2757( .A (n218), .B (n219), .C (n90), .Y (n2765) );
  AO21x1_ASAP7_75t_R   g2758( .A1 (n1300), .A2 (n217), .B (n2765), .Y (n2766) );
  INVx1_ASAP7_75t_R    g2759( .A (n2766), .Y (n2767) );
  AND2x2_ASAP7_75t_R   g2760( .A (n64), .B (n84), .Y (n2768) );
  AND2x2_ASAP7_75t_R   g2761( .A (n2767), .B (n2768), .Y (y1118) );
  OA211x2_ASAP7_75t_R  g2762( .A1 (n2710), .A2 (n1885), .B (n2736), .C (n84), .Y (y1119) );
  AND2x2_ASAP7_75t_R   g2763( .A (n2414), .B (n2768), .Y (y1120) );
  AND2x2_ASAP7_75t_R   g2764( .A (n84), .B (n64), .Y (n2772) );
  NAND2x1_ASAP7_75t_R  g2765( .A (x1), .B (n863), .Y (n2773) );
  AND2x2_ASAP7_75t_R   g2766( .A (n2772), .B (n2773), .Y (y1121) );
  AO21x1_ASAP7_75t_R   g2767( .A1 (n17), .A2 (x0), .B (n392), .Y (n2775) );
  INVx1_ASAP7_75t_R    g2768( .A (n2775), .Y (n2776) );
  OR3x1_ASAP7_75t_R    g2769( .A (n315), .B (y2079), .C (x3), .Y (n2777) );
  INVx1_ASAP7_75t_R    g2770( .A (n2777), .Y (n2778) );
  AO21x1_ASAP7_75t_R   g2771( .A1 (n391), .A2 (n2776), .B (n2778), .Y (n2779) );
  AO21x1_ASAP7_75t_R   g2772( .A1 (x0), .A2 (x4), .B (n2779), .Y (y1122) );
  AND3x1_ASAP7_75t_R   g2773( .A (n17), .B (n12), .C (x1), .Y (n2781) );
  NOR2x1_ASAP7_75t_R   g2774( .A (n1536), .B (n2756), .Y (n2782) );
  AO21x1_ASAP7_75t_R   g2775( .A1 (x2), .A2 (n2781), .B (n2782), .Y (y1123) );
  NAND2x1_ASAP7_75t_R  g2776( .A (n2038), .B (n64), .Y (n2784) );
  OAI21x1_ASAP7_75t_R  g2777( .A1 (n12), .A2 (n2784), .B (x3), .Y (n2785) );
  OA21x2_ASAP7_75t_R   g2778( .A1 (x3), .A2 (n2784), .B (n2785), .Y (y1124) );
  AO21x1_ASAP7_75t_R   g2779( .A1 (x3), .A2 (x2), .B (n16), .Y (n2787) );
  AND2x2_ASAP7_75t_R   g2780( .A (n2787), .B (x0), .Y (n2788) );
  AND3x1_ASAP7_75t_R   g2781( .A (n16), .B (x3), .C (x2), .Y (n2789) );
  INVx1_ASAP7_75t_R    g2782( .A (n2789), .Y (n2790) );
  OA21x2_ASAP7_75t_R   g2783( .A1 (n2788), .A2 (n81), .B (n2790), .Y (y1125) );
  AND3x1_ASAP7_75t_R   g2784( .A (x0), .B (x3), .C (x2), .Y (n2792) );
  INVx1_ASAP7_75t_R    g2785( .A (n2792), .Y (n2793) );
  AO21x1_ASAP7_75t_R   g2786( .A1 (n2793), .A2 (n1572), .B (n16), .Y (n2794) );
  NAND2x1_ASAP7_75t_R  g2787( .A (n806), .B (n2794), .Y (y1126) );
  OA21x2_ASAP7_75t_R   g2788( .A1 (n382), .A2 (n363), .B (n1997), .Y (n2796) );
  OR3x1_ASAP7_75t_R    g2789( .A (n145), .B (x5), .C (x4), .Y (n2797) );
  OA21x2_ASAP7_75t_R   g2790( .A1 (n2796), .A2 (x0), .B (n2797), .Y (y1127) );
  AO21x1_ASAP7_75t_R   g2791( .A1 (n16), .A2 (n2137), .B (n2147), .Y (y1128) );
  OR3x1_ASAP7_75t_R    g2792( .A (n2583), .B (n826), .C (x3), .Y (n2800) );
  AO21x1_ASAP7_75t_R   g2793( .A1 (n827), .A2 (n1301), .B (n17), .Y (n2801) );
  AND2x2_ASAP7_75t_R   g2794( .A (n2800), .B (n2801), .Y (n2802) );
  NOR2x1_ASAP7_75t_R   g2795( .A (n1032), .B (n2802), .Y (y1129) );
  AO21x1_ASAP7_75t_R   g2796( .A1 (n72), .A2 (n137), .B (n90), .Y (n2804) );
  NAND2x1_ASAP7_75t_R  g2797( .A (n2804), .B (n2794), .Y (y1130) );
  AO21x1_ASAP7_75t_R   g2798( .A1 (n2060), .A2 (x1), .B (n58), .Y (y1131) );
  AO21x1_ASAP7_75t_R   g2799( .A1 (n125), .A2 (x2), .B (n1656), .Y (n2807) );
  AND2x2_ASAP7_75t_R   g2800( .A (n805), .B (n2807), .Y (y1132) );
  AO21x1_ASAP7_75t_R   g2801( .A1 (n90), .A2 (n211), .B (n2546), .Y (n2809) );
  AO21x1_ASAP7_75t_R   g2802( .A1 (n12), .A2 (x3), .B (x2), .Y (n2810) );
  NOR2x1_ASAP7_75t_R   g2803( .A (x1), .B (n2810), .Y (n2811) );
  AO21x1_ASAP7_75t_R   g2804( .A1 (n2809), .A2 (x0), .B (n2811), .Y (y1133) );
  AND3x1_ASAP7_75t_R   g2805( .A (n63), .B (n64), .C (n17), .Y (n2813) );
  INVx1_ASAP7_75t_R    g2806( .A (n2813), .Y (n2814) );
  AND3x1_ASAP7_75t_R   g2807( .A (n2814), .B (n1671), .C (x0), .Y (y1135) );
  AO21x1_ASAP7_75t_R   g2808( .A1 (n1391), .A2 (n2407), .B (y2079), .Y (y1136) );
  AO21x1_ASAP7_75t_R   g2809( .A1 (n378), .A2 (y2079), .B (x0), .Y (y1137) );
  AO21x1_ASAP7_75t_R   g2810( .A1 (n12), .A2 (n15), .B (n13), .Y (n2818) );
  AO21x1_ASAP7_75t_R   g2811( .A1 (n970), .A2 (n2818), .B (n730), .Y (y1138) );
  AO21x1_ASAP7_75t_R   g2812( .A1 (n12), .A2 (n15), .B (x1), .Y (n2820) );
  AO21x1_ASAP7_75t_R   g2813( .A1 (n2820), .A2 (n2158), .B (y2093), .Y (y1139) );
  OR3x1_ASAP7_75t_R    g2814( .A (y2093), .B (n262), .C (n1649), .Y (y1140) );
  AO21x1_ASAP7_75t_R   g2815( .A1 (y2079), .A2 (n797), .B (n754), .Y (y1141) );
  OR3x1_ASAP7_75t_R    g2816( .A (n2147), .B (y2196), .C (n61), .Y (y1142) );
  NAND2x1_ASAP7_75t_R  g2817( .A (n12), .B (n878), .Y (n2825) );
  XOR2x2_ASAP7_75t_R   g2818( .A (n1676), .B (n2825), .Y (y1143) );
  AND3x1_ASAP7_75t_R   g2819( .A (y2079), .B (x1), .C (x0), .Y (y2022) );
  AO21x1_ASAP7_75t_R   g2820( .A1 (n12), .A2 (n16), .B (y2022), .Y (n2828) );
  AO21x1_ASAP7_75t_R   g2821( .A1 (n2828), .A2 (n15), .B (n2156), .Y (y1144) );
  AND2x2_ASAP7_75t_R   g2822( .A (n221), .B (n164), .Y (n2830) );
  AO21x1_ASAP7_75t_R   g2823( .A1 (x2), .A2 (n1668), .B (n2830), .Y (y1145) );
  AO21x1_ASAP7_75t_R   g2824( .A1 (y2079), .A2 (x0), .B (n51), .Y (n2832) );
  NAND2x1_ASAP7_75t_R  g2825( .A (n51), .B (y3852), .Y (n2833) );
  OA21x2_ASAP7_75t_R   g2826( .A1 (n2147), .A2 (n2832), .B (n2833), .Y (y1146) );
  OA21x2_ASAP7_75t_R   g2827( .A1 (n65), .A2 (n1510), .B (n2516), .Y (y1147) );
  OR3x1_ASAP7_75t_R    g2828( .A (n43), .B (y2079), .C (n103), .Y (n2836) );
  AND2x2_ASAP7_75t_R   g2829( .A (n2836), .B (n244), .Y (y1148) );
  AND3x1_ASAP7_75t_R   g2830( .A (n1870), .B (n1640), .C (n244), .Y (y1149) );
  INVx1_ASAP7_75t_R    g2831( .A (n1521), .Y (n2839) );
  NOR2x1_ASAP7_75t_R   g2832( .A (n1462), .B (n2839), .Y (y1150) );
  AND3x1_ASAP7_75t_R   g2833( .A (x1), .B (x3), .C (x2), .Y (n2841) );
  OR3x1_ASAP7_75t_R    g2834( .A (n2841), .B (n81), .C (x0), .Y (y1151) );
  INVx1_ASAP7_75t_R    g2835( .A (n2027), .Y (n2843) );
  AO21x1_ASAP7_75t_R   g2836( .A1 (n2843), .A2 (n16), .B (n143), .Y (y1152) );
  OA21x2_ASAP7_75t_R   g2837( .A1 (n1644), .A2 (n2508), .B (n1246), .Y (y1153) );
  AO21x1_ASAP7_75t_R   g2838( .A1 (n1530), .A2 (n497), .B (n109), .Y (y1154) );
  AO21x1_ASAP7_75t_R   g2839( .A1 (n12), .A2 (n17), .B (x2), .Y (n2847) );
  AO21x1_ASAP7_75t_R   g2840( .A1 (n16), .A2 (n15), .B (x3), .Y (n2848) );
  AND2x2_ASAP7_75t_R   g2841( .A (n2848), .B (x0), .Y (n2849) );
  AO21x1_ASAP7_75t_R   g2842( .A1 (n2847), .A2 (x1), .B (n2849), .Y (y1155) );
  OA21x2_ASAP7_75t_R   g2843( .A1 (n1644), .A2 (n2508), .B (n1870), .Y (y1156) );
  OA21x2_ASAP7_75t_R   g2844( .A1 (n1437), .A2 (x1), .B (n1332), .Y (y1157) );
  NOR2x1_ASAP7_75t_R   g2845( .A (x1), .B (n751), .Y (n2853) );
  OR3x1_ASAP7_75t_R    g2846( .A (n2853), .B (n856), .C (n2169), .Y (y1158) );
  AO32x1_ASAP7_75t_R   g2847( .A1 (n1954), .A2 (n913), .A3 (n15), .B1 (x2), .B2 (y873), .Y (y1159) );
  OA211x2_ASAP7_75t_R  g2848( .A1 (n2140), .A2 (y2196), .B (n2509), .C (n219), .Y (y1160) );
  OA21x2_ASAP7_75t_R   g2849( .A1 (n771), .A2 (n2508), .B (n90), .Y (y1161) );
  AO32x1_ASAP7_75t_R   g2850( .A1 (n15), .A2 (n144), .A3 (n913), .B1 (x2), .B2 (y873), .Y (y1162) );
  AO21x1_ASAP7_75t_R   g2851( .A1 (n97), .A2 (y1356), .B (n2126), .Y (y1163) );
  NAND2x1_ASAP7_75t_R  g2852( .A (n565), .B (n219), .Y (n2860) );
  AO33x2_ASAP7_75t_R   g2853( .A1 (n219), .A2 (n565), .A3 (x2), .B1 (n2860), .B2 (n15), .B3 (n913), .Y (y1164) );
  AND2x2_ASAP7_75t_R   g2854( .A (n2404), .B (n2117), .Y (y1165) );
  AND3x1_ASAP7_75t_R   g2855( .A (n97), .B (n64), .C (x0), .Y (y1207) );
  AO21x1_ASAP7_75t_R   g2856( .A1 (n128), .A2 (n481), .B (y1207), .Y (y1166) );
  INVx1_ASAP7_75t_R    g2857( .A (n175), .Y (n2865) );
  AO21x1_ASAP7_75t_R   g2858( .A1 (n2508), .A2 (x1), .B (n2865), .Y (y1167) );
  AO21x1_ASAP7_75t_R   g2859( .A1 (n1305), .A2 (n271), .B (n262), .Y (y1168) );
  NAND2x1_ASAP7_75t_R  g2860( .A (x3), .B (n185), .Y (n2868) );
  AO32x1_ASAP7_75t_R   g2861( .A1 (n228), .A2 (n2868), .A3 (n2258), .B1 (x2), .B2 (n1682), .Y (y1169) );
  AO21x1_ASAP7_75t_R   g2862( .A1 (n765), .A2 (n51), .B (n2441), .Y (y1170) );
  AO21x1_ASAP7_75t_R   g2863( .A1 (x2), .A2 (x0), .B (n16), .Y (n2871) );
  AO21x1_ASAP7_75t_R   g2864( .A1 (n15), .A2 (n12), .B (x1), .Y (n2872) );
  NAND2x1_ASAP7_75t_R  g2865( .A (n2871), .B (n2872), .Y (n2873) );
  INVx1_ASAP7_75t_R    g2866( .A (n2873), .Y (y1171) );
  AND3x1_ASAP7_75t_R   g2867( .A (n64), .B (n219), .C (n2810), .Y (y1172) );
  AO21x1_ASAP7_75t_R   g2868( .A1 (x1), .A2 (x2), .B (n12), .Y (n2876) );
  NAND2x1_ASAP7_75t_R  g2869( .A (n2876), .B (n1457), .Y (n2877) );
  AO21x1_ASAP7_75t_R   g2870( .A1 (n12), .A2 (x2), .B (n17), .Y (n2878) );
  AO21x1_ASAP7_75t_R   g2871( .A1 (y9), .A2 (n2679), .B (n2878), .Y (n2879) );
  INVx1_ASAP7_75t_R    g2872( .A (n2879), .Y (n2880) );
  AO21x1_ASAP7_75t_R   g2873( .A1 (n17), .A2 (n2877), .B (n2880), .Y (y1173) );
  AND3x1_ASAP7_75t_R   g2874( .A (n72), .B (n90), .C (n219), .Y (n2882) );
  AO21x1_ASAP7_75t_R   g2875( .A1 (n17), .A2 (x2), .B (n227), .Y (n2883) );
  XOR2x2_ASAP7_75t_R   g2876( .A (n2882), .B (n2883), .Y (y1174) );
  OR3x1_ASAP7_75t_R    g2877( .A (n51), .B (y2079), .C (x0), .Y (n2885) );
  AO21x1_ASAP7_75t_R   g2878( .A1 (n15), .A2 (n16), .B (y2079), .Y (n2886) );
  AO21x1_ASAP7_75t_R   g2879( .A1 (n2886), .A2 (x0), .B (n13), .Y (n2887) );
  AO21x1_ASAP7_75t_R   g2880( .A1 (n2885), .A2 (n2887), .B (n1587), .Y (y1175) );
  INVx1_ASAP7_75t_R    g2881( .A (n1295), .Y (n2889) );
  OA33x2_ASAP7_75t_R   g2882( .A1 (x2), .A2 (n2889), .A3 (n43), .B1 (n111), .B2 (n15), .B3 (n2565), .Y (y1176) );
  AO21x1_ASAP7_75t_R   g2883( .A1 (n12), .A2 (x1), .B (n17), .Y (n2891) );
  AO21x1_ASAP7_75t_R   g2884( .A1 (n242), .A2 (n14), .B (n2891), .Y (n2892) );
  INVx1_ASAP7_75t_R    g2885( .A (n2892), .Y (n2893) );
  AO21x1_ASAP7_75t_R   g2886( .A1 (n17), .A2 (n1676), .B (n2893), .Y (y1177) );
  AND3x1_ASAP7_75t_R   g2887( .A (n700), .B (n757), .C (n63), .Y (n2895) );
  OR2x4_ASAP7_75t_R    g2888( .A (x0), .B (n2895), .Y (n2896) );
  AND3x1_ASAP7_75t_R   g2889( .A (n58), .B (n16), .C (n15), .Y (n2897) );
  INVx1_ASAP7_75t_R    g2890( .A (n2897), .Y (n2898) );
  AND2x2_ASAP7_75t_R   g2891( .A (n2896), .B (n2898), .Y (y1178) );
  OR3x1_ASAP7_75t_R    g2892( .A (n43), .B (n17), .C (n103), .Y (n2900) );
  OA21x2_ASAP7_75t_R   g2893( .A1 (n145), .A2 (n1301), .B (n2900), .Y (y1179) );
  AO21x1_ASAP7_75t_R   g2894( .A1 (n1295), .A2 (n1296), .B (x2), .Y (n2902) );
  INVx1_ASAP7_75t_R    g2895( .A (n2902), .Y (n2903) );
  AO21x1_ASAP7_75t_R   g2896( .A1 (n17), .A2 (x1), .B (n12), .Y (n2904) );
  INVx1_ASAP7_75t_R    g2897( .A (n2904), .Y (n2905) );
  AO21x1_ASAP7_75t_R   g2898( .A1 (n72), .A2 (x1), .B (n133), .Y (n2906) );
  OA21x2_ASAP7_75t_R   g2899( .A1 (n2903), .A2 (n2905), .B (n2906), .Y (y1180) );
  AO21x1_ASAP7_75t_R   g2900( .A1 (n17), .A2 (x0), .B (n43), .Y (n2908) );
  AO21x1_ASAP7_75t_R   g2901( .A1 (n1301), .A2 (n2908), .B (n2544), .Y (y1181) );
  OR3x1_ASAP7_75t_R    g2902( .A (n13), .B (n17), .C (n12), .Y (n2910) );
  NAND2x1_ASAP7_75t_R  g2903( .A (n17), .B (n703), .Y (n2911) );
  AND3x1_ASAP7_75t_R   g2904( .A (n2910), .B (n2911), .C (n67), .Y (y1182) );
  OR3x1_ASAP7_75t_R    g2905( .A (n241), .B (y2079), .C (x1), .Y (n2913) );
  INVx1_ASAP7_75t_R    g2906( .A (n2913), .Y (n2914) );
  AO21x1_ASAP7_75t_R   g2907( .A1 (n1340), .A2 (n497), .B (n12), .Y (n2915) );
  OA21x2_ASAP7_75t_R   g2908( .A1 (n2914), .A2 (n2699), .B (n2915), .Y (y1183) );
  INVx1_ASAP7_75t_R    g2909( .A (n210), .Y (n2917) );
  OR3x1_ASAP7_75t_R    g2910( .A (n163), .B (n164), .C (n12), .Y (n2918) );
  AOI22x1_ASAP7_75t_R  g2911( .A1 (n2917), .A2 (n191), .B1 (n210), .B2 (n2918), .Y (y1184) );
  AND2x2_ASAP7_75t_R   g2912( .A (n1455), .B (n706), .Y (y1185) );
  INVx1_ASAP7_75t_R    g2913( .A (n883), .Y (n2921) );
  AO21x1_ASAP7_75t_R   g2914( .A1 (n17), .A2 (n15), .B (y863), .Y (n2922) );
  AO21x1_ASAP7_75t_R   g2915( .A1 (n2921), .A2 (n12), .B (n2922), .Y (n2923) );
  NAND2x1_ASAP7_75t_R  g2916( .A (n2923), .B (n2273), .Y (n2924) );
  INVx1_ASAP7_75t_R    g2917( .A (n2924), .Y (y1186) );
  AO21x1_ASAP7_75t_R   g2918( .A1 (y863), .A2 (x2), .B (y2079), .Y (y1187) );
  AND3x1_ASAP7_75t_R   g2919( .A (n14), .B (n67), .C (y2079), .Y (n2927) );
  NOR2x1_ASAP7_75t_R   g2920( .A (n481), .B (n2927), .Y (y1188) );
  AND3x1_ASAP7_75t_R   g2921( .A (x2), .B (x1), .C (x0), .Y (y1214) );
  AO21x1_ASAP7_75t_R   g2922( .A1 (y0), .A2 (y2079), .B (y1214), .Y (y1189) );
  AO21x1_ASAP7_75t_R   g2923( .A1 (n103), .A2 (x0), .B (y2079), .Y (n2931) );
  AND2x2_ASAP7_75t_R   g2924( .A (n187), .B (n2931), .Y (y1190) );
  AO21x1_ASAP7_75t_R   g2925( .A1 (y9), .A2 (y2079), .B (n2169), .Y (y1191) );
  AO21x1_ASAP7_75t_R   g2926( .A1 (y2079), .A2 (y25), .B (n2441), .Y (y1192) );
  AO21x1_ASAP7_75t_R   g2927( .A1 (x2), .A2 (n143), .B (n2347), .Y (y1193) );
  AND2x2_ASAP7_75t_R   g2928( .A (y1193), .B (n52), .Y (y1194) );
  AND2x2_ASAP7_75t_R   g2929( .A (n244), .B (n2172), .Y (y1195) );
  AND3x1_ASAP7_75t_R   g2930( .A (n1870), .B (n244), .C (n97), .Y (y1196) );
  AO21x1_ASAP7_75t_R   g2931( .A1 (n497), .A2 (n276), .B (n1339), .Y (y1197) );
  OR3x1_ASAP7_75t_R    g2932( .A (n58), .B (n16), .C (x4), .Y (n2940) );
  AND3x1_ASAP7_75t_R   g2933( .A (n1246), .B (n2940), .C (n299), .Y (y1198) );
  OA21x2_ASAP7_75t_R   g2934( .A1 (n993), .A2 (n2511), .B (n2182), .Y (y1200) );
  AO21x1_ASAP7_75t_R   g2935( .A1 (n497), .A2 (n276), .B (n801), .Y (y1202) );
  AO21x1_ASAP7_75t_R   g2936( .A1 (n174), .A2 (y2079), .B (n262), .Y (y1203) );
  AO21x1_ASAP7_75t_R   g2937( .A1 (n12), .A2 (n705), .B (y1207), .Y (y1204) );
  AO21x1_ASAP7_75t_R   g2938( .A1 (x1), .A2 (n276), .B (n856), .Y (y1205) );
  AND3x1_ASAP7_75t_R   g2939( .A (n97), .B (n244), .C (n851), .Y (y1206) );
  AO21x1_ASAP7_75t_R   g2940( .A1 (n16), .A2 (n242), .B (n1208), .Y (n2948) );
  NOR2x1_ASAP7_75t_R   g2941( .A (n1646), .B (n2948), .Y (y1208) );
  OA21x2_ASAP7_75t_R   g2942( .A1 (x0), .A2 (n1173), .B (n1001), .Y (y1209) );
  AO21x1_ASAP7_75t_R   g2943( .A1 (n173), .A2 (n856), .B (n262), .Y (y1210) );
  AO21x1_ASAP7_75t_R   g2944( .A1 (n16), .A2 (n15), .B (x5), .Y (n2952) );
  INVx1_ASAP7_75t_R    g2945( .A (n2952), .Y (n2953) );
  OA21x2_ASAP7_75t_R   g2946( .A1 (n2953), .A2 (n2315), .B (n2675), .Y (y1211) );
  OA21x2_ASAP7_75t_R   g2947( .A1 (n94), .A2 (n13), .B (x0), .Y (y1212) );
  AND3x1_ASAP7_75t_R   g2948( .A (n64), .B (n219), .C (n2136), .Y (y1213) );
  AO21x1_ASAP7_75t_R   g2949( .A1 (n103), .A2 (x0), .B (n17), .Y (n2957) );
  OA21x2_ASAP7_75t_R   g2950( .A1 (n1693), .A2 (x3), .B (n2957), .Y (y1215) );
  INVx1_ASAP7_75t_R    g2951( .A (n244), .Y (n2959) );
  OR3x1_ASAP7_75t_R    g2952( .A (n2959), .B (x5), .C (x1), .Y (n2960) );
  AND2x2_ASAP7_75t_R   g2953( .A (n2960), .B (y3852), .Y (y1216) );
  AO21x1_ASAP7_75t_R   g2954( .A1 (n998), .A2 (n15), .B (n2496), .Y (y1217) );
  OR3x1_ASAP7_75t_R    g2955( .A (n45), .B (y2079), .C (x4), .Y (n2963) );
  INVx1_ASAP7_75t_R    g2956( .A (n2963), .Y (n2964) );
  AND3x1_ASAP7_75t_R   g2957( .A (x2), .B (x3), .C (x5), .Y (n2965) );
  INVx1_ASAP7_75t_R    g2958( .A (n2965), .Y (n2966) );
  OA21x2_ASAP7_75t_R   g2959( .A1 (n2964), .A2 (n211), .B (n2966), .Y (y1218) );
  AND3x1_ASAP7_75t_R   g2960( .A (n2490), .B (n2069), .C (n64), .Y (y1219) );
  NOR2x1_ASAP7_75t_R   g2961( .A (x2), .B (n1997), .Y (n2969) );
  INVx1_ASAP7_75t_R    g2962( .A (n2969), .Y (n2970) );
  AO21x1_ASAP7_75t_R   g2963( .A1 (n17), .A2 (n15), .B (y2079), .Y (n2971) );
  AO21x1_ASAP7_75t_R   g2964( .A1 (n77), .A2 (n22), .B (n2971), .Y (y1267) );
  AND2x2_ASAP7_75t_R   g2965( .A (n2970), .B (y1267), .Y (y1220) );
  OR3x1_ASAP7_75t_R    g2966( .A (n529), .B (n29), .C (n1093), .Y (n2974) );
  AND2x2_ASAP7_75t_R   g2967( .A (n2974), .B (n602), .Y (y1221) );
  AO21x1_ASAP7_75t_R   g2968( .A1 (n17), .A2 (n56), .B (n813), .Y (y1222) );
  NAND2x1_ASAP7_75t_R  g2969( .A (n740), .B (n746), .Y (n2977) );
  OA21x2_ASAP7_75t_R   g2970( .A1 (x1), .A2 (n2977), .B (n2612), .Y (y1223) );
  OR3x1_ASAP7_75t_R    g2971( .A (n325), .B (y2079), .C (x2), .Y (n2979) );
  AO21x1_ASAP7_75t_R   g2972( .A1 (x4), .A2 (x3), .B (x2), .Y (n2980) );
  AO21x1_ASAP7_75t_R   g2973( .A1 (y2079), .A2 (n2980), .B (n347), .Y (n2981) );
  NOR2x1_ASAP7_75t_R   g2974( .A (x2), .B (n2049), .Y (n2982) );
  AO21x1_ASAP7_75t_R   g2975( .A1 (n2979), .A2 (n2981), .B (n2982), .Y (y1224) );
  AO21x1_ASAP7_75t_R   g2976( .A1 (n299), .A2 (n310), .B (x3), .Y (n2984) );
  OA21x2_ASAP7_75t_R   g2977( .A1 (n291), .A2 (y1281), .B (n2984), .Y (y1225) );
  NAND2x1_ASAP7_75t_R  g2978( .A (x4), .B (n1242), .Y (n2986) );
  OR3x1_ASAP7_75t_R    g2979( .A (n1380), .B (n227), .C (x4), .Y (n2987) );
  AND2x2_ASAP7_75t_R   g2980( .A (n2986), .B (n2987), .Y (y1226) );
  AND3x1_ASAP7_75t_R   g2981( .A (n22), .B (x3), .C (x2), .Y (n2989) );
  AO21x1_ASAP7_75t_R   g2982( .A1 (x5), .A2 (n2989), .B (n529), .Y (n2990) );
  AO21x1_ASAP7_75t_R   g2983( .A1 (n45), .A2 (n28), .B (n2990), .Y (y1227) );
  AO21x1_ASAP7_75t_R   g2984( .A1 (n290), .A2 (n360), .B (n12), .Y (n2992) );
  INVx1_ASAP7_75t_R    g2985( .A (n2992), .Y (n2993) );
  AND3x1_ASAP7_75t_R   g2986( .A (n17), .B (x4), .C (x0), .Y (n2994) );
  NOR2x1_ASAP7_75t_R   g2987( .A (x5), .B (n2994), .Y (n2995) );
  AO21x1_ASAP7_75t_R   g2988( .A1 (n2993), .A2 (x5), .B (n2995), .Y (y1228) );
  AND3x1_ASAP7_75t_R   g2989( .A (n137), .B (n72), .C (x5), .Y (n2997) );
  AO21x1_ASAP7_75t_R   g2990( .A1 (x3), .A2 (x2), .B (n22), .Y (n2998) );
  NOR2x1_ASAP7_75t_R   g2991( .A (x2), .B (x4), .Y (n2999) );
  INVx1_ASAP7_75t_R    g2992( .A (n2999), .Y (n3000) );
  AO21x1_ASAP7_75t_R   g2993( .A1 (n15), .A2 (x3), .B (y2079), .Y (n3001) );
  AO21x1_ASAP7_75t_R   g2994( .A1 (n3000), .A2 (n17), .B (n3001), .Y (n3002) );
  OA21x2_ASAP7_75t_R   g2995( .A1 (n2997), .A2 (n2998), .B (n3002), .Y (y1229) );
  AO21x1_ASAP7_75t_R   g2996( .A1 (n12), .A2 (n17), .B (n368), .Y (n3004) );
  INVx1_ASAP7_75t_R    g2997( .A (n3004), .Y (n3005) );
  AO21x1_ASAP7_75t_R   g2998( .A1 (n583), .A2 (n17), .B (n650), .Y (n3006) );
  INVx1_ASAP7_75t_R    g2999( .A (n3006), .Y (n3007) );
  AO21x1_ASAP7_75t_R   g3000( .A1 (x4), .A2 (n3005), .B (n3007), .Y (y1230) );
  AND3x1_ASAP7_75t_R   g3001( .A (n22), .B (x5), .C (x3), .Y (n3009) );
  AO21x1_ASAP7_75t_R   g3002( .A1 (n3005), .A2 (x4), .B (n3009), .Y (y1231) );
  AO21x1_ASAP7_75t_R   g3003( .A1 (x5), .A2 (x4), .B (x2), .Y (n3011) );
  AND3x1_ASAP7_75t_R   g3004( .A (x2), .B (x5), .C (x4), .Y (n3012) );
  INVx1_ASAP7_75t_R    g3005( .A (n3012), .Y (n3013) );
  AO21x1_ASAP7_75t_R   g3006( .A1 (y2079), .A2 (n22), .B (n17), .Y (n3014) );
  AO32x1_ASAP7_75t_R   g3007( .A1 (n3011), .A2 (n3013), .A3 (n3014), .B1 (y3293), .B2 (n164), .Y (y1232) );
  INVx1_ASAP7_75t_R    g3008( .A (n2470), .Y (n3016) );
  OA21x2_ASAP7_75t_R   g3009( .A1 (x1), .A2 (n3016), .B (n2605), .Y (y1233) );
  OR3x1_ASAP7_75t_R    g3010( .A (n2050), .B (n2051), .C (x2), .Y (n3018) );
  AO21x1_ASAP7_75t_R   g3011( .A1 (n660), .A2 (n406), .B (n15), .Y (n3019) );
  AND2x2_ASAP7_75t_R   g3012( .A (n3018), .B (n3019), .Y (y1234) );
  AO21x1_ASAP7_75t_R   g3013( .A1 (n1271), .A2 (n22), .B (n1078), .Y (n3021) );
  AND2x2_ASAP7_75t_R   g3014( .A (n3021), .B (n1272), .Y (y1235) );
  AO21x1_ASAP7_75t_R   g3015( .A1 (n15), .A2 (n17), .B (y2079), .Y (n3023) );
  AO21x1_ASAP7_75t_R   g3016( .A1 (x2), .A2 (x3), .B (x4), .Y (n3024) );
  INVx1_ASAP7_75t_R    g3017( .A (n3024), .Y (n3025) );
  NAND2x1_ASAP7_75t_R  g3018( .A (n3023), .B (n3025), .Y (n3026) );
  AND2x2_ASAP7_75t_R   g3019( .A (x2), .B (x4), .Y (n3027) );
  INVx1_ASAP7_75t_R    g3020( .A (n3027), .Y (n3028) );
  AO21x1_ASAP7_75t_R   g3021( .A1 (n15), .A2 (n22), .B (y2079), .Y (n3029) );
  AO21x1_ASAP7_75t_R   g3022( .A1 (n3028), .A2 (n17), .B (n3029), .Y (n3030) );
  AND3x1_ASAP7_75t_R   g3023( .A (n3026), .B (n3030), .C (n1265), .Y (y1236) );
  AND2x2_ASAP7_75t_R   g3024( .A (n738), .B (n827), .Y (y1237) );
  INVx1_ASAP7_75t_R    g3025( .A (n2810), .Y (n3033) );
  AO21x1_ASAP7_75t_R   g3026( .A1 (n12), .A2 (x2), .B (n16), .Y (n3034) );
  INVx1_ASAP7_75t_R    g3027( .A (n3034), .Y (n3035) );
  AO21x1_ASAP7_75t_R   g3028( .A1 (n125), .A2 (n16), .B (n2810), .Y (n3036) );
  OA21x2_ASAP7_75t_R   g3029( .A1 (n3033), .A2 (n3035), .B (n3036), .Y (y1238) );
  AO21x1_ASAP7_75t_R   g3030( .A1 (n29), .A2 (y9), .B (n529), .Y (y1239) );
  AO21x1_ASAP7_75t_R   g3031( .A1 (n139), .A2 (n22), .B (n325), .Y (n3039) );
  AO21x1_ASAP7_75t_R   g3032( .A1 (x4), .A2 (x3), .B (n12), .Y (n3040) );
  NAND2x1_ASAP7_75t_R  g3033( .A (x5), .B (n3040), .Y (y3176) );
  OA21x2_ASAP7_75t_R   g3034( .A1 (x5), .A2 (n3039), .B (y3176), .Y (y1240) );
  AO21x1_ASAP7_75t_R   g3035( .A1 (n15), .A2 (n17), .B (n12), .Y (n3043) );
  NAND2x1_ASAP7_75t_R  g3036( .A (n3043), .B (n165), .Y (y1241) );
  AO21x1_ASAP7_75t_R   g3037( .A1 (n16), .A2 (n12), .B (n392), .Y (n3045) );
  INVx1_ASAP7_75t_R    g3038( .A (n3045), .Y (y1242) );
  NAND2x1_ASAP7_75t_R  g3039( .A (n17), .B (n1775), .Y (n3047) );
  AND2x2_ASAP7_75t_R   g3040( .A (n3047), .B (y168), .Y (y1243) );
  NAND2x1_ASAP7_75t_R  g3041( .A (n12), .B (n523), .Y (n3049) );
  INVx1_ASAP7_75t_R    g3042( .A (n727), .Y (n3050) );
  AO21x1_ASAP7_75t_R   g3043( .A1 (n3049), .A2 (y3293), .B (n3050), .Y (y1244) );
  OR3x1_ASAP7_75t_R    g3044( .A (n1016), .B (n529), .C (n527), .Y (y1245) );
  AND2x2_ASAP7_75t_R   g3045( .A (n3049), .B (y3293), .Y (y1246) );
  AO21x1_ASAP7_75t_R   g3046( .A1 (x0), .A2 (n17), .B (n28), .Y (n3054) );
  INVx1_ASAP7_75t_R    g3047( .A (n3054), .Y (n3055) );
  AO21x1_ASAP7_75t_R   g3048( .A1 (n28), .A2 (n3005), .B (n3055), .Y (y1247) );
  NAND2x1_ASAP7_75t_R  g3049( .A (n2008), .B (n781), .Y (n3057) );
  AND2x2_ASAP7_75t_R   g3050( .A (n3057), .B (y3293), .Y (y1248) );
  NOR2x1_ASAP7_75t_R   g3051( .A (y2466), .B (n900), .Y (y1249) );
  AND3x1_ASAP7_75t_R   g3052( .A (y103), .B (n934), .C (n17), .Y (n3060) );
  OR3x1_ASAP7_75t_R    g3053( .A (n392), .B (n17), .C (n12), .Y (n3061) );
  INVx1_ASAP7_75t_R    g3054( .A (n3061), .Y (n3062) );
  OR3x1_ASAP7_75t_R    g3055( .A (n3060), .B (n3062), .C (n418), .Y (y1250) );
  AND3x1_ASAP7_75t_R   g3056( .A (n137), .B (n72), .C (n16), .Y (n3064) );
  INVx1_ASAP7_75t_R    g3057( .A (n3043), .Y (n3065) );
  OA21x2_ASAP7_75t_R   g3058( .A1 (n3064), .A2 (n3065), .B (n90), .Y (y1251) );
  AO32x1_ASAP7_75t_R   g3059( .A1 (y2079), .A2 (n244), .A3 (n16), .B1 (x1), .B2 (n707), .Y (y1252) );
  AND2x2_ASAP7_75t_R   g3060( .A (y3758), .B (y9), .Y (y1253) );
  AO21x1_ASAP7_75t_R   g3061( .A1 (n388), .A2 (n28), .B (n15), .Y (n3069) );
  INVx1_ASAP7_75t_R    g3062( .A (n3069), .Y (n3070) );
  AO21x1_ASAP7_75t_R   g3063( .A1 (n3070), .A2 (x3), .B (n81), .Y (y1254) );
  AO21x1_ASAP7_75t_R   g3064( .A1 (n12), .A2 (x3), .B (x4), .Y (n3072) );
  AND2x2_ASAP7_75t_R   g3065( .A (n3072), .B (y2079), .Y (n3073) );
  AO21x1_ASAP7_75t_R   g3066( .A1 (n22), .A2 (n397), .B (n3073), .Y (y1255) );
  AO21x1_ASAP7_75t_R   g3067( .A1 (n378), .A2 (x5), .B (n2051), .Y (y1260) );
  AND2x2_ASAP7_75t_R   g3068( .A (y1260), .B (x0), .Y (y1256) );
  OR3x1_ASAP7_75t_R    g3069( .A (n139), .B (y2079), .C (n403), .Y (n3077) );
  NAND2x1_ASAP7_75t_R  g3070( .A (n388), .B (n3077), .Y (y1257) );
  AO21x1_ASAP7_75t_R   g3071( .A1 (n16), .A2 (n1646), .B (n1503), .Y (y1258) );
  AND3x1_ASAP7_75t_R   g3072( .A (n22), .B (x3), .C (x0), .Y (n3080) );
  OR3x1_ASAP7_75t_R    g3073( .A (n1775), .B (n3080), .C (n638), .Y (y1259) );
  AO21x1_ASAP7_75t_R   g3074( .A1 (n29), .A2 (n84), .B (n1775), .Y (y1261) );
  AO21x1_ASAP7_75t_R   g3075( .A1 (n15), .A2 (x3), .B (x5), .Y (n3083) );
  NOR2x1_ASAP7_75t_R   g3076( .A (n3027), .B (n3083), .Y (y1262) );
  INVx1_ASAP7_75t_R    g3077( .A (n3072), .Y (n3085) );
  AO21x1_ASAP7_75t_R   g3078( .A1 (n3085), .A2 (n352), .B (n529), .Y (y1263) );
  AO21x1_ASAP7_75t_R   g3079( .A1 (n29), .A2 (n84), .B (n529), .Y (y1264) );
  NAND2x1_ASAP7_75t_R  g3080( .A (x5), .B (n3072), .Y (y1343) );
  OR3x1_ASAP7_75t_R    g3081( .A (x0), .B (x3), .C (x5), .Y (n3089) );
  AND2x2_ASAP7_75t_R   g3082( .A (y1343), .B (n3089), .Y (y1265) );
  INVx1_ASAP7_75t_R    g3083( .A (n978), .Y (n3091) );
  AND3x1_ASAP7_75t_R   g3084( .A (n2182), .B (n2701), .C (n3091), .Y (y1266) );
  AO21x1_ASAP7_75t_R   g3085( .A1 (n455), .A2 (x0), .B (n363), .Y (n3093) );
  AND2x2_ASAP7_75t_R   g3086( .A (n3093), .B (n1114), .Y (y1268) );
  AND3x1_ASAP7_75t_R   g3087( .A (n84), .B (n22), .C (x5), .Y (n3095) );
  AO21x1_ASAP7_75t_R   g3088( .A1 (y2079), .A2 (n2645), .B (n3095), .Y (y1269) );
  AO21x1_ASAP7_75t_R   g3089( .A1 (x2), .A2 (x5), .B (n17), .Y (n3097) );
  AO32x1_ASAP7_75t_R   g3090( .A1 (n3028), .A2 (n3097), .A3 (n388), .B1 (n529), .B2 (n1062), .Y (y1270) );
  INVx1_ASAP7_75t_R    g3091( .A (n639), .Y (n3099) );
  AO21x1_ASAP7_75t_R   g3092( .A1 (n29), .A2 (n84), .B (n3099), .Y (y1271) );
  AND3x1_ASAP7_75t_R   g3093( .A (n556), .B (n290), .C (n360), .Y (n3101) );
  AO21x1_ASAP7_75t_R   g3094( .A1 (n556), .A2 (x0), .B (n3101), .Y (y1272) );
  AO21x1_ASAP7_75t_R   g3095( .A1 (n63), .A2 (n752), .B (n754), .Y (y1273) );
  OA21x2_ASAP7_75t_R   g3096( .A1 (n397), .A2 (n403), .B (n556), .Y (y1274) );
  INVx1_ASAP7_75t_R    g3097( .A (n351), .Y (n3105) );
  OA21x2_ASAP7_75t_R   g3098( .A1 (n3105), .A2 (n1319), .B (n357), .Y (y1275) );
  NOR2x1_ASAP7_75t_R   g3099( .A (n139), .B (n388), .Y (n3107) );
  AO21x1_ASAP7_75t_R   g3100( .A1 (n84), .A2 (n29), .B (n3107), .Y (y1276) );
  OR3x1_ASAP7_75t_R    g3101( .A (n325), .B (n12), .C (x5), .Y (n3109) );
  AND3x1_ASAP7_75t_R   g3102( .A (n3109), .B (y672), .C (y3377), .Y (y1277) );
  AO21x1_ASAP7_75t_R   g3103( .A1 (n63), .A2 (y2079), .B (n143), .Y (y1278) );
  AND2x2_ASAP7_75t_R   g3104( .A (n125), .B (y2079), .Y (n3112) );
  OA22x2_ASAP7_75t_R   g3105( .A1 (n421), .A2 (n1851), .B1 (n3112), .B2 (n22), .Y (y1279) );
  NAND2x1_ASAP7_75t_R  g3106( .A (n3072), .B (n388), .Y (y1777) );
  AND2x2_ASAP7_75t_R   g3107( .A (y1777), .B (n645), .Y (y1280) );
  INVx1_ASAP7_75t_R    g3108( .A (n2645), .Y (n3116) );
  NAND2x1_ASAP7_75t_R  g3109( .A (n510), .B (n3116), .Y (n3117) );
  AND3x1_ASAP7_75t_R   g3110( .A (x3), .B (x4), .C (x5), .Y (n3118) );
  INVx1_ASAP7_75t_R    g3111( .A (n3118), .Y (n3119) );
  AND2x2_ASAP7_75t_R   g3112( .A (n3117), .B (n3119), .Y (y1282) );
  AO21x1_ASAP7_75t_R   g3113( .A1 (n12), .A2 (x4), .B (n145), .Y (n3121) );
  OA21x2_ASAP7_75t_R   g3114( .A1 (n421), .A2 (n3121), .B (n556), .Y (y1284) );
  AO21x1_ASAP7_75t_R   g3115( .A1 (n15), .A2 (y2079), .B (x4), .Y (n3123) );
  INVx1_ASAP7_75t_R    g3116( .A (n3123), .Y (n3124) );
  AO21x1_ASAP7_75t_R   g3117( .A1 (n3124), .A2 (n1838), .B (n529), .Y (y1285) );
  AO21x1_ASAP7_75t_R   g3118( .A1 (n352), .A2 (n51), .B (y1201), .Y (y1286) );
  OR3x1_ASAP7_75t_R    g3119( .A (n529), .B (n29), .C (n45), .Y (y1287) );
  AO21x1_ASAP7_75t_R   g3120( .A1 (n17), .A2 (x0), .B (n22), .Y (n3128) );
  NOR2x1_ASAP7_75t_R   g3121( .A (x5), .B (n3128), .Y (n3129) );
  AO21x1_ASAP7_75t_R   g3122( .A1 (n84), .A2 (n29), .B (n3129), .Y (y1288) );
  AO21x1_ASAP7_75t_R   g3123( .A1 (n16), .A2 (n572), .B (n957), .Y (y1289) );
  AND3x1_ASAP7_75t_R   g3124( .A (y2079), .B (x2), .C (x3), .Y (n3132) );
  AO21x1_ASAP7_75t_R   g3125( .A1 (n17), .A2 (n15), .B (n3132), .Y (n3133) );
  AO21x1_ASAP7_75t_R   g3126( .A1 (n137), .A2 (n72), .B (x4), .Y (n3134) );
  INVx1_ASAP7_75t_R    g3127( .A (n3134), .Y (n3135) );
  AO21x1_ASAP7_75t_R   g3128( .A1 (n3133), .A2 (x4), .B (n3135), .Y (y1290) );
  AND2x2_ASAP7_75t_R   g3129( .A (n2971), .B (n2998), .Y (y1291) );
  OR3x1_ASAP7_75t_R    g3130( .A (n529), .B (n29), .C (n1158), .Y (n3138) );
  OR3x1_ASAP7_75t_R    g3131( .A (y2466), .B (n17), .C (x0), .Y (n3139) );
  AND2x2_ASAP7_75t_R   g3132( .A (n3138), .B (n3139), .Y (y1292) );
  AND3x1_ASAP7_75t_R   g3133( .A (n2999), .B (n17), .C (x5), .Y (n3141) );
  AO21x1_ASAP7_75t_R   g3134( .A1 (y2079), .A2 (n1572), .B (n3141), .Y (y1293) );
  AO21x1_ASAP7_75t_R   g3135( .A1 (x3), .A2 (x4), .B (x2), .Y (n3143) );
  INVx1_ASAP7_75t_R    g3136( .A (n3143), .Y (n3144) );
  AND2x2_ASAP7_75t_R   g3137( .A (n406), .B (x2), .Y (n3145) );
  AO21x1_ASAP7_75t_R   g3138( .A1 (n1997), .A2 (n3144), .B (n3145), .Y (y1294) );
  NAND2x1_ASAP7_75t_R  g3139( .A (x3), .B (n430), .Y (n3147) );
  OR3x1_ASAP7_75t_R    g3140( .A (x0), .B (x5), .C (x4), .Y (n3148) );
  INVx1_ASAP7_75t_R    g3141( .A (n3148), .Y (n3149) );
  AO21x1_ASAP7_75t_R   g3142( .A1 (n3147), .A2 (y3293), .B (n3149), .Y (y1295) );
  AND2x2_ASAP7_75t_R   g3143( .A (n3147), .B (y3293), .Y (y1296) );
  AND2x2_ASAP7_75t_R   g3144( .A (y3758), .B (n84), .Y (y1297) );
  AND2x2_ASAP7_75t_R   g3145( .A (n1176), .B (y2079), .Y (y1298) );
  NAND2x1_ASAP7_75t_R  g3146( .A (n697), .B (n310), .Y (y1299) );
  AO32x1_ASAP7_75t_R   g3147( .A1 (y2079), .A2 (n436), .A3 (n1853), .B1 (x5), .B2 (n1176), .Y (y1301) );
  INVx1_ASAP7_75t_R    g3148( .A (y1116), .Y (n3156) );
  AO21x1_ASAP7_75t_R   g3149( .A1 (n16), .A2 (x5), .B (n276), .Y (n3157) );
  AND2x2_ASAP7_75t_R   g3150( .A (n3157), .B (n64), .Y (n3158) );
  AO21x1_ASAP7_75t_R   g3151( .A1 (n3156), .A2 (y2079), .B (n3158), .Y (y1302) );
  AO21x1_ASAP7_75t_R   g3152( .A1 (n12), .A2 (x3), .B (x5), .Y (n3160) );
  OA21x2_ASAP7_75t_R   g3153( .A1 (n537), .A2 (n3160), .B (y1343), .Y (y1303) );
  AND2x2_ASAP7_75t_R   g3154( .A (y117), .B (n469), .Y (y1304) );
  AO21x1_ASAP7_75t_R   g3155( .A1 (n14), .A2 (x3), .B (n235), .Y (n3163) );
  INVx1_ASAP7_75t_R    g3156( .A (n3163), .Y (n3164) );
  AND3x1_ASAP7_75t_R   g3157( .A (n3164), .B (n52), .C (x0), .Y (y1305) );
  OR3x1_ASAP7_75t_R    g3158( .A (n139), .B (x5), .C (x4), .Y (n3166) );
  AND2x2_ASAP7_75t_R   g3159( .A (n3166), .B (y1281), .Y (y1306) );
  AO21x1_ASAP7_75t_R   g3160( .A1 (n17), .A2 (x2), .B (n392), .Y (n3168) );
  INVx1_ASAP7_75t_R    g3161( .A (n3168), .Y (n3169) );
  OR3x1_ASAP7_75t_R    g3162( .A (x2), .B (x5), .C (x4), .Y (n3170) );
  AO21x1_ASAP7_75t_R   g3163( .A1 (n3169), .A2 (n3170), .B (n297), .Y (y1307) );
  AND2x2_ASAP7_75t_R   g3164( .A (n1997), .B (x0), .Y (n3172) );
  NAND2x1_ASAP7_75t_R  g3165( .A (n12), .B (n641), .Y (n3173) );
  INVx1_ASAP7_75t_R    g3166( .A (n3173), .Y (n3174) );
  AO21x1_ASAP7_75t_R   g3167( .A1 (n3119), .A2 (n3172), .B (n3174), .Y (y1309) );
  NAND2x1_ASAP7_75t_R  g3168( .A (x4), .B (n1106), .Y (n3176) );
  OA21x2_ASAP7_75t_R   g3169( .A1 (x4), .A2 (n530), .B (n3176), .Y (y1310) );
  AO21x1_ASAP7_75t_R   g3170( .A1 (n1387), .A2 (n1060), .B (n1266), .Y (y1311) );
  NAND2x1_ASAP7_75t_R  g3171( .A (n1106), .B (n310), .Y (y1997) );
  AND2x2_ASAP7_75t_R   g3172( .A (y1997), .B (n451), .Y (y1312) );
  AO21x1_ASAP7_75t_R   g3173( .A1 (n22), .A2 (x2), .B (x3), .Y (n3181) );
  INVx1_ASAP7_75t_R    g3174( .A (n3181), .Y (n3182) );
  AO21x1_ASAP7_75t_R   g3175( .A1 (n15), .A2 (x4), .B (y2079), .Y (n3183) );
  AO21x1_ASAP7_75t_R   g3176( .A1 (x2), .A2 (x5), .B (x3), .Y (n3184) );
  AO21x1_ASAP7_75t_R   g3177( .A1 (n3124), .A2 (n3184), .B (n529), .Y (n3185) );
  AO21x1_ASAP7_75t_R   g3178( .A1 (n3182), .A2 (n3183), .B (n3185), .Y (y1313) );
  AND3x1_ASAP7_75t_R   g3179( .A (n2940), .B (y9), .C (n556), .Y (y1314) );
  AO21x1_ASAP7_75t_R   g3180( .A1 (n2814), .A2 (n1671), .B (x0), .Y (y1315) );
  AND3x1_ASAP7_75t_R   g3181( .A (n22), .B (n17), .C (x0), .Y (n3189) );
  AO21x1_ASAP7_75t_R   g3182( .A1 (n348), .A2 (n363), .B (n3189), .Y (y1316) );
  AO21x1_ASAP7_75t_R   g3183( .A1 (x0), .A2 (x5), .B (n17), .Y (n3191) );
  AND3x1_ASAP7_75t_R   g3184( .A (n17), .B (x5), .C (x0), .Y (n3192) );
  AO21x1_ASAP7_75t_R   g3185( .A1 (y2079), .A2 (x3), .B (n3192), .Y (n3193) );
  AO21x1_ASAP7_75t_R   g3186( .A1 (n22), .A2 (n3191), .B (n3193), .Y (y1317) );
  AO21x1_ASAP7_75t_R   g3187( .A1 (n388), .A2 (n28), .B (n90), .Y (n3195) );
  AND2x2_ASAP7_75t_R   g3188( .A (n3195), .B (y104), .Y (y1318) );
  INVx1_ASAP7_75t_R    g3189( .A (n1007), .Y (n3197) );
  OR3x1_ASAP7_75t_R    g3190( .A (n43), .B (y2079), .C (n22), .Y (n3198) );
  OA21x2_ASAP7_75t_R   g3191( .A1 (n3197), .A2 (n58), .B (n3198), .Y (y1319) );
  AO21x1_ASAP7_75t_R   g3192( .A1 (n740), .A2 (n43), .B (y742), .Y (y1320) );
  AO21x1_ASAP7_75t_R   g3193( .A1 (x2), .A2 (y2079), .B (n173), .Y (n3201) );
  AO32x1_ASAP7_75t_R   g3194( .A1 (y2079), .A2 (n187), .A3 (n3201), .B1 (x5), .B2 (y2393), .Y (y1321) );
  INVx1_ASAP7_75t_R    g3195( .A (n299), .Y (n3203) );
  OR3x1_ASAP7_75t_R    g3196( .A (n3203), .B (x5), .C (x1), .Y (n3204) );
  AND2x2_ASAP7_75t_R   g3197( .A (n3204), .B (y1281), .Y (y1322) );
  AO21x1_ASAP7_75t_R   g3198( .A1 (n596), .A2 (y2079), .B (n914), .Y (y1323) );
  AO21x1_ASAP7_75t_R   g3199( .A1 (n17), .A2 (x5), .B (x4), .Y (n3207) );
  NAND2x1_ASAP7_75t_R  g3200( .A (n3207), .B (n290), .Y (n3208) );
  OR3x1_ASAP7_75t_R    g3201( .A (n337), .B (y2079), .C (n15), .Y (n3209) );
  OA21x2_ASAP7_75t_R   g3202( .A1 (n3208), .A2 (x2), .B (n3209), .Y (y1324) );
  AND3x1_ASAP7_75t_R   g3203( .A (n369), .B (n370), .C (x0), .Y (n3211) );
  INVx1_ASAP7_75t_R    g3204( .A (n3211), .Y (n3212) );
  AO21x1_ASAP7_75t_R   g3205( .A1 (y3852), .A2 (n17), .B (n718), .Y (n3213) );
  AND3x1_ASAP7_75t_R   g3206( .A (n3212), .B (n3213), .C (y3852), .Y (y1325) );
  INVx1_ASAP7_75t_R    g3207( .A (n589), .Y (n3215) );
  OA211x2_ASAP7_75t_R  g3208( .A1 (n1851), .A2 (n231), .B (n3215), .C (n556), .Y (y1326) );
  AND2x2_ASAP7_75t_R   g3209( .A (n443), .B (n1125), .Y (y1327) );
  AND3x1_ASAP7_75t_R   g3210( .A (x5), .B (x4), .C (x3), .Y (n3218) );
  NOR2x1_ASAP7_75t_R   g3211( .A (n12), .B (n3218), .Y (y1328) );
  AND2x2_ASAP7_75t_R   g3212( .A (y1300), .B (n3215), .Y (y1329) );
  NAND2x1_ASAP7_75t_R  g3213( .A (n976), .B (n388), .Y (y1330) );
  AO21x1_ASAP7_75t_R   g3214( .A1 (x1), .A2 (x4), .B (n12), .Y (n3222) );
  NAND2x1_ASAP7_75t_R  g3215( .A (y2079), .B (n3222), .Y (n3223) );
  INVx1_ASAP7_75t_R    g3216( .A (n3223), .Y (n3224) );
  AO21x1_ASAP7_75t_R   g3217( .A1 (n22), .A2 (n1093), .B (n3224), .Y (y1331) );
  AO21x1_ASAP7_75t_R   g3218( .A1 (y2079), .A2 (n899), .B (n905), .Y (y1332) );
  AND3x1_ASAP7_75t_R   g3219( .A (n290), .B (n360), .C (n15), .Y (n3227) );
  INVx1_ASAP7_75t_R    g3220( .A (n3209), .Y (n3228) );
  NOR2x1_ASAP7_75t_R   g3221( .A (n3227), .B (n3228), .Y (y1333) );
  AO21x1_ASAP7_75t_R   g3222( .A1 (y2079), .A2 (n90), .B (n914), .Y (y2832) );
  AND2x2_ASAP7_75t_R   g3223( .A (y2832), .B (n451), .Y (y1334) );
  AND3x1_ASAP7_75t_R   g3224( .A (n43), .B (n15), .C (x5), .Y (n3232) );
  INVx1_ASAP7_75t_R    g3225( .A (n3232), .Y (y1335) );
  AND3x1_ASAP7_75t_R   g3226( .A (y2079), .B (x3), .C (x0), .Y (n3234) );
  AO21x1_ASAP7_75t_R   g3227( .A1 (n17), .A2 (n22), .B (n3234), .Y (y1336) );
  NAND2x1_ASAP7_75t_R  g3228( .A (n2199), .B (n794), .Y (y1337) );
  AO21x1_ASAP7_75t_R   g3229( .A1 (y2079), .A2 (x4), .B (n15), .Y (n3237) );
  AO21x1_ASAP7_75t_R   g3230( .A1 (n388), .A2 (n17), .B (x2), .Y (n3238) );
  OA21x2_ASAP7_75t_R   g3231( .A1 (n3237), .A2 (n3009), .B (n3238), .Y (y1338) );
  AND2x2_ASAP7_75t_R   g3232( .A (y1300), .B (n700), .Y (y1339) );
  AO21x1_ASAP7_75t_R   g3233( .A1 (n1246), .A2 (n750), .B (n495), .Y (n3241) );
  AND2x2_ASAP7_75t_R   g3234( .A (n3241), .B (n244), .Y (y1340) );
  AND2x2_ASAP7_75t_R   g3235( .A (n488), .B (n22), .Y (n3243) );
  OA21x2_ASAP7_75t_R   g3236( .A1 (n3243), .A2 (y2196), .B (n1026), .Y (y1341) );
  AND3x1_ASAP7_75t_R   g3237( .A (n1863), .B (y1281), .C (n466), .Y (y1342) );
  AND2x2_ASAP7_75t_R   g3238( .A (n2661), .B (n2172), .Y (y1344) );
  NOR2x1_ASAP7_75t_R   g3239( .A (n16), .B (n614), .Y (n3247) );
  AO21x1_ASAP7_75t_R   g3240( .A1 (n22), .A2 (n1093), .B (n3247), .Y (y1345) );
  NOR2x1_ASAP7_75t_R   g3241( .A (x5), .B (x0), .Y (n3249) );
  AND2x2_ASAP7_75t_R   g3242( .A (x5), .B (x0), .Y (n3250) );
  AND3x1_ASAP7_75t_R   g3243( .A (n3250), .B (n17), .C (n22), .Y (n3251) );
  AO21x1_ASAP7_75t_R   g3244( .A1 (n377), .A2 (n3249), .B (n3251), .Y (y1346) );
  AO21x1_ASAP7_75t_R   g3245( .A1 (y3852), .A2 (n1163), .B (n437), .Y (n3253) );
  AND2x2_ASAP7_75t_R   g3246( .A (n1863), .B (n3253), .Y (y1347) );
  AO21x1_ASAP7_75t_R   g3247( .A1 (n914), .A2 (x5), .B (n1907), .Y (y1348) );
  NAND2x1_ASAP7_75t_R  g3248( .A (n337), .B (n352), .Y (n3256) );
  INVx1_ASAP7_75t_R    g3249( .A (n3256), .Y (n3257) );
  AO21x1_ASAP7_75t_R   g3250( .A1 (y2079), .A2 (n2645), .B (n3257), .Y (y1349) );
  AND2x2_ASAP7_75t_R   g3251( .A (y3852), .B (n436), .Y (n3259) );
  AO21x1_ASAP7_75t_R   g3252( .A1 (n28), .A2 (n3259), .B (n503), .Y (y1350) );
  NAND2x1_ASAP7_75t_R  g3253( .A (x4), .B (n3160), .Y (n3261) );
  OA21x2_ASAP7_75t_R   g3254( .A1 (n628), .A2 (n1851), .B (n3261), .Y (y1351) );
  AND3x1_ASAP7_75t_R   g3255( .A (n15), .B (n17), .C (x4), .Y (n3263) );
  AO21x1_ASAP7_75t_R   g3256( .A1 (n15), .A2 (n17), .B (n392), .Y (n3264) );
  NOR2x1_ASAP7_75t_R   g3257( .A (n959), .B (n3264), .Y (n3265) );
  AO21x1_ASAP7_75t_R   g3258( .A1 (x5), .A2 (n3263), .B (n3265), .Y (y1352) );
  AO21x1_ASAP7_75t_R   g3259( .A1 (n22), .A2 (x0), .B (x3), .Y (n3267) );
  INVx1_ASAP7_75t_R    g3260( .A (n3267), .Y (n3268) );
  NOR2x1_ASAP7_75t_R   g3261( .A (n12), .B (n671), .Y (n3269) );
  OA21x2_ASAP7_75t_R   g3262( .A1 (n3268), .A2 (n3269), .B (y1281), .Y (y1353) );
  NAND2x1_ASAP7_75t_R  g3263( .A (n45), .B (n28), .Y (n3271) );
  INVx1_ASAP7_75t_R    g3264( .A (n3271), .Y (n3272) );
  AO21x1_ASAP7_75t_R   g3265( .A1 (y3758), .A2 (x2), .B (n3272), .Y (y1354) );
  OR3x1_ASAP7_75t_R    g3266( .A (n58), .B (x4), .C (x3), .Y (n3274) );
  AO21x1_ASAP7_75t_R   g3267( .A1 (n12), .A2 (x3), .B (n518), .Y (n3275) );
  INVx1_ASAP7_75t_R    g3268( .A (n3275), .Y (n3276) );
  AND2x2_ASAP7_75t_R   g3269( .A (n3274), .B (n3276), .Y (y1355) );
  AO21x1_ASAP7_75t_R   g3270( .A1 (y2079), .A2 (x2), .B (n45), .Y (n3278) );
  AND3x1_ASAP7_75t_R   g3271( .A (n22), .B (x5), .C (x2), .Y (n3279) );
  AO21x1_ASAP7_75t_R   g3272( .A1 (n3278), .A2 (x4), .B (n3279), .Y (y1357) );
  AO21x1_ASAP7_75t_R   g3273( .A1 (n466), .A2 (n58), .B (n1071), .Y (y1358) );
  AO21x1_ASAP7_75t_R   g3274( .A1 (x3), .A2 (x2), .B (x4), .Y (n3282) );
  NAND2x1_ASAP7_75t_R  g3275( .A (x5), .B (n3282), .Y (y1359) );
  AO21x1_ASAP7_75t_R   g3276( .A1 (n17), .A2 (x5), .B (n22), .Y (n3284) );
  AO21x1_ASAP7_75t_R   g3277( .A1 (y2079), .A2 (x3), .B (n15), .Y (n3285) );
  NAND2x1_ASAP7_75t_R  g3278( .A (n15), .B (n3284), .Y (n3286) );
  OA21x2_ASAP7_75t_R   g3279( .A1 (n3284), .A2 (n3285), .B (n3286), .Y (y1360) );
  AO21x1_ASAP7_75t_R   g3280( .A1 (n84), .A2 (n125), .B (n103), .Y (n3288) );
  AO21x1_ASAP7_75t_R   g3281( .A1 (n15), .A2 (n626), .B (n3288), .Y (y1361) );
  AO21x1_ASAP7_75t_R   g3282( .A1 (n299), .A2 (n310), .B (n17), .Y (n3290) );
  INVx1_ASAP7_75t_R    g3283( .A (n3290), .Y (n3291) );
  NAND2x1_ASAP7_75t_R  g3284( .A (y2079), .B (n3291), .Y (n3292) );
  AND2x2_ASAP7_75t_R   g3285( .A (n3292), .B (y1281), .Y (y1362) );
  AND3x1_ASAP7_75t_R   g3286( .A (n15), .B (n17), .C (x5), .Y (n3294) );
  NAND2x1_ASAP7_75t_R  g3287( .A (x4), .B (n3294), .Y (n3295) );
  INVx1_ASAP7_75t_R    g3288( .A (n3295), .Y (n3296) );
  AO21x1_ASAP7_75t_R   g3289( .A1 (x4), .A2 (x5), .B (n15), .Y (n3297) );
  INVx1_ASAP7_75t_R    g3290( .A (n3297), .Y (n3298) );
  OR3x1_ASAP7_75t_R    g3291( .A (n3296), .B (n3298), .C (n628), .Y (y1363) );
  OA21x2_ASAP7_75t_R   g3292( .A1 (n316), .A2 (n537), .B (y1281), .Y (y1364) );
  INVx1_ASAP7_75t_R    g3293( .A (n366), .Y (n3301) );
  NAND2x1_ASAP7_75t_R  g3294( .A (x2), .B (n3301), .Y (n3302) );
  AND2x2_ASAP7_75t_R   g3295( .A (n3302), .B (n72), .Y (y1365) );
  INVx1_ASAP7_75t_R    g3296( .A (n835), .Y (n3304) );
  OA21x2_ASAP7_75t_R   g3297( .A1 (n3304), .A2 (n988), .B (n2296), .Y (n3305) );
  AO21x1_ASAP7_75t_R   g3298( .A1 (y2079), .A2 (x0), .B (n3305), .Y (y1366) );
  AND3x1_ASAP7_75t_R   g3299( .A (n1838), .B (n64), .C (n63), .Y (n3307) );
  AND3x1_ASAP7_75t_R   g3300( .A (n152), .B (n153), .C (x0), .Y (y3968) );
  AO21x1_ASAP7_75t_R   g3301( .A1 (n12), .A2 (n3307), .B (y3968), .Y (y1367) );
  AND3x1_ASAP7_75t_R   g3302( .A (n15), .B (x4), .C (x3), .Y (n3310) );
  NOR2x1_ASAP7_75t_R   g3303( .A (n347), .B (n3310), .Y (n3311) );
  AND3x1_ASAP7_75t_R   g3304( .A (n347), .B (n15), .C (x5), .Y (n3312) );
  AO21x1_ASAP7_75t_R   g3305( .A1 (n3311), .A2 (y2079), .B (n3312), .Y (y1368) );
  AND3x1_ASAP7_75t_R   g3306( .A (y194), .B (n546), .C (n463), .Y (y1369) );
  AND3x1_ASAP7_75t_R   g3307( .A (x4), .B (x3), .C (x2), .Y (n3315) );
  INVx1_ASAP7_75t_R    g3308( .A (n3282), .Y (n3316) );
  NOR2x1_ASAP7_75t_R   g3309( .A (n3315), .B (n3316), .Y (n3317) );
  NAND2x1_ASAP7_75t_R  g3310( .A (n81), .B (n388), .Y (n3318) );
  OA21x2_ASAP7_75t_R   g3311( .A1 (n3317), .A2 (y2079), .B (n3318), .Y (y1370) );
  AND3x1_ASAP7_75t_R   g3312( .A (y9), .B (y1894), .C (y3293), .Y (y1371) );
  OR3x1_ASAP7_75t_R    g3313( .A (n530), .B (n2458), .C (x4), .Y (n3321) );
  AND2x2_ASAP7_75t_R   g3314( .A (n3321), .B (n3176), .Y (y1372) );
  OR3x1_ASAP7_75t_R    g3315( .A (n143), .B (x2), .C (x3), .Y (n3323) );
  NAND2x1_ASAP7_75t_R  g3316( .A (n2684), .B (n3323), .Y (y1373) );
  AO21x1_ASAP7_75t_R   g3317( .A1 (n12), .A2 (x4), .B (x3), .Y (n3325) );
  AO21x1_ASAP7_75t_R   g3318( .A1 (n310), .A2 (x5), .B (n3325), .Y (n3326) );
  AO21x1_ASAP7_75t_R   g3319( .A1 (n17), .A2 (x0), .B (y2079), .Y (n3327) );
  AO21x1_ASAP7_75t_R   g3320( .A1 (n84), .A2 (n22), .B (n3327), .Y (y2727) );
  AND2x2_ASAP7_75t_R   g3321( .A (n3326), .B (y2727), .Y (y1374) );
  INVx1_ASAP7_75t_R    g3322( .A (n2551), .Y (y1375) );
  OR3x1_ASAP7_75t_R    g3323( .A (n529), .B (n29), .C (n437), .Y (n3331) );
  AND2x2_ASAP7_75t_R   g3324( .A (n3331), .B (n2016), .Y (y1376) );
  AND3x1_ASAP7_75t_R   g3325( .A (n15), .B (x3), .C (x4), .Y (n3333) );
  INVx1_ASAP7_75t_R    g3326( .A (n3333), .Y (n3334) );
  AND2x2_ASAP7_75t_R   g3327( .A (n3209), .B (n3334), .Y (y1377) );
  AO21x1_ASAP7_75t_R   g3328( .A1 (n231), .A2 (n22), .B (x0), .Y (n3336) );
  AND3x1_ASAP7_75t_R   g3329( .A (n445), .B (n3336), .C (n556), .Y (y1379) );
  AO21x1_ASAP7_75t_R   g3330( .A1 (n22), .A2 (x5), .B (n17), .Y (n3338) );
  AO22x1_ASAP7_75t_R   g3331( .A1 (n3183), .A2 (x3), .B1 (n3338), .B2 (x2), .Y (y1380) );
  AND2x2_ASAP7_75t_R   g3332( .A (n3331), .B (x0), .Y (y1381) );
  AND2x2_ASAP7_75t_R   g3333( .A (n660), .B (n661), .Y (n3341) );
  NOR2x1_ASAP7_75t_R   g3334( .A (x5), .B (n3341), .Y (n3342) );
  AO21x1_ASAP7_75t_R   g3335( .A1 (n3191), .A2 (n474), .B (n3342), .Y (y1382) );
  INVx1_ASAP7_75t_R    g3336( .A (n3080), .Y (n3344) );
  AO21x1_ASAP7_75t_R   g3337( .A1 (n3344), .A2 (n299), .B (x5), .Y (n3345) );
  AND2x2_ASAP7_75t_R   g3338( .A (n3345), .B (y1281), .Y (y1383) );
  AND3x1_ASAP7_75t_R   g3339( .A (n1370), .B (n718), .C (y3852), .Y (y1384) );
  AND3x1_ASAP7_75t_R   g3340( .A (y1359), .B (n455), .C (n1572), .Y (y1385) );
  AO21x1_ASAP7_75t_R   g3341( .A1 (y2079), .A2 (x1), .B (n15), .Y (n3349) );
  AO21x1_ASAP7_75t_R   g3342( .A1 (n497), .A2 (x0), .B (n3349), .Y (n3350) );
  OA21x2_ASAP7_75t_R   g3343( .A1 (n1815), .A2 (x2), .B (n3350), .Y (y1386) );
  AO21x1_ASAP7_75t_R   g3344( .A1 (n22), .A2 (x0), .B (n1907), .Y (y1387) );
  AND2x2_ASAP7_75t_R   g3345( .A (n3013), .B (n72), .Y (y1388) );
  INVx1_ASAP7_75t_R    g3346( .A (n959), .Y (n3354) );
  AND3x1_ASAP7_75t_R   g3347( .A (n3354), .B (y3293), .C (x0), .Y (y1389) );
  OR3x1_ASAP7_75t_R    g3348( .A (n1380), .B (n227), .C (x2), .Y (n3356) );
  NAND2x1_ASAP7_75t_R  g3349( .A (n2258), .B (n3356), .Y (y1390) );
  AND2x2_ASAP7_75t_R   g3350( .A (y3758), .B (x0), .Y (y1391) );
  AO21x1_ASAP7_75t_R   g3351( .A1 (n22), .A2 (x5), .B (n15), .Y (n3359) );
  AO21x1_ASAP7_75t_R   g3352( .A1 (y2079), .A2 (x4), .B (n17), .Y (n3360) );
  NOR2x1_ASAP7_75t_R   g3353( .A (n3359), .B (n3360), .Y (n3361) );
  NOR2x1_ASAP7_75t_R   g3354( .A (n81), .B (n3361), .Y (y1392) );
  NAND2x1_ASAP7_75t_R  g3355( .A (x5), .B (n1306), .Y (y1393) );
  AO21x1_ASAP7_75t_R   g3356( .A1 (n3182), .A2 (n1265), .B (n293), .Y (y1394) );
  INVx1_ASAP7_75t_R    g3357( .A (n490), .Y (n3365) );
  OR3x1_ASAP7_75t_R    g3358( .A (x0), .B (x1), .C (x4), .Y (n3366) );
  AND2x2_ASAP7_75t_R   g3359( .A (n3366), .B (y2079), .Y (n3367) );
  AO21x1_ASAP7_75t_R   g3360( .A1 (n3365), .A2 (n970), .B (n3367), .Y (y1395) );
  AO21x1_ASAP7_75t_R   g3361( .A1 (n17), .A2 (y2079), .B (n12), .Y (n3369) );
  AO21x1_ASAP7_75t_R   g3362( .A1 (n12), .A2 (n17), .B (n22), .Y (n3370) );
  NAND2x1_ASAP7_75t_R  g3363( .A (n3369), .B (n3370), .Y (n3371) );
  OR3x1_ASAP7_75t_R    g3364( .A (n671), .B (n22), .C (n12), .Y (n3372) );
  AND3x1_ASAP7_75t_R   g3365( .A (n3371), .B (n3372), .C (n369), .Y (y1396) );
  AO21x1_ASAP7_75t_R   g3366( .A1 (n15), .A2 (x4), .B (x3), .Y (n3374) );
  INVx1_ASAP7_75t_R    g3367( .A (n3374), .Y (n3375) );
  AO21x1_ASAP7_75t_R   g3368( .A1 (x3), .A2 (x4), .B (x5), .Y (n3376) );
  AO21x1_ASAP7_75t_R   g3369( .A1 (n17), .A2 (x4), .B (x2), .Y (n3377) );
  AO21x1_ASAP7_75t_R   g3370( .A1 (n3028), .A2 (n3377), .B (y2079), .Y (y3276) );
  OA21x2_ASAP7_75t_R   g3371( .A1 (n3375), .A2 (n3376), .B (y3276), .Y (y1397) );
  NAND2x1_ASAP7_75t_R  g3372( .A (x5), .B (n490), .Y (n3380) );
  AND2x2_ASAP7_75t_R   g3373( .A (n3380), .B (n2940), .Y (y1398) );
  AO21x1_ASAP7_75t_R   g3374( .A1 (x1), .A2 (n58), .B (n43), .Y (n3382) );
  AO21x1_ASAP7_75t_R   g3375( .A1 (n22), .A2 (n3382), .B (n529), .Y (y1399) );
  INVx1_ASAP7_75t_R    g3376( .A (n3128), .Y (n3384) );
  NAND2x1_ASAP7_75t_R  g3377( .A (x5), .B (n3384), .Y (y1903) );
  AND3x1_ASAP7_75t_R   g3378( .A (n17), .B (n22), .C (x0), .Y (n3386) );
  INVx1_ASAP7_75t_R    g3379( .A (n3386), .Y (n3387) );
  AND2x2_ASAP7_75t_R   g3380( .A (y1903), .B (n3387), .Y (y2144) );
  OA21x2_ASAP7_75t_R   g3381( .A1 (x5), .A2 (n3384), .B (y2144), .Y (y1400) );
  NOR2x1_ASAP7_75t_R   g3382( .A (n316), .B (n310), .Y (n3390) );
  INVx1_ASAP7_75t_R    g3383( .A (n3390), .Y (n3391) );
  NAND2x1_ASAP7_75t_R  g3384( .A (n639), .B (n310), .Y (n3392) );
  AND2x2_ASAP7_75t_R   g3385( .A (n3391), .B (n3392), .Y (y1401) );
  AO21x1_ASAP7_75t_R   g3386( .A1 (n1923), .A2 (n90), .B (y2079), .Y (n3394) );
  AO21x1_ASAP7_75t_R   g3387( .A1 (n466), .A2 (n436), .B (x0), .Y (n3395) );
  AND2x2_ASAP7_75t_R   g3388( .A (n3394), .B (n3395), .Y (y1402) );
  OA21x2_ASAP7_75t_R   g3389( .A1 (n1819), .A2 (n478), .B (n546), .Y (y1403) );
  AO21x1_ASAP7_75t_R   g3390( .A1 (x0), .A2 (y2079), .B (n290), .Y (n3398) );
  INVx1_ASAP7_75t_R    g3391( .A (n3398), .Y (n3399) );
  AO21x1_ASAP7_75t_R   g3392( .A1 (n556), .A2 (n351), .B (n3399), .Y (y1404) );
  AO21x1_ASAP7_75t_R   g3393( .A1 (y2079), .A2 (x4), .B (n905), .Y (y2878) );
  AND2x2_ASAP7_75t_R   g3394( .A (y2878), .B (n1385), .Y (y1405) );
  AO21x1_ASAP7_75t_R   g3395( .A1 (y855), .A2 (n228), .B (y2079), .Y (y1406) );
  AO21x1_ASAP7_75t_R   g3396( .A1 (n22), .A2 (x0), .B (n16), .Y (n3404) );
  AND3x1_ASAP7_75t_R   g3397( .A (n90), .B (n3404), .C (y2079), .Y (n3405) );
  INVx1_ASAP7_75t_R    g3398( .A (n3405), .Y (n3406) );
  AND2x2_ASAP7_75t_R   g3399( .A (y1393), .B (n3406), .Y (y1407) );
  AO21x1_ASAP7_75t_R   g3400( .A1 (x1), .A2 (n22), .B (n604), .Y (y1845) );
  AND2x2_ASAP7_75t_R   g3401( .A (y1845), .B (n546), .Y (y1408) );
  AND2x2_ASAP7_75t_R   g3402( .A (n2940), .B (n556), .Y (n3410) );
  AND2x2_ASAP7_75t_R   g3403( .A (n1410), .B (n3410), .Y (y1409) );
  NAND2x1_ASAP7_75t_R  g3404( .A (y2079), .B (n948), .Y (n3412) );
  AND2x2_ASAP7_75t_R   g3405( .A (y1393), .B (n3412), .Y (y1410) );
  INVx1_ASAP7_75t_R    g3406( .A (n334), .Y (n3414) );
  OA21x2_ASAP7_75t_R   g3407( .A1 (n315), .A2 (x3), .B (y2079), .Y (n3415) );
  AO21x1_ASAP7_75t_R   g3408( .A1 (n3414), .A2 (x5), .B (n3415), .Y (y1411) );
  NOR2x1_ASAP7_75t_R   g3409( .A (x5), .B (n315), .Y (n3417) );
  OA21x2_ASAP7_75t_R   g3410( .A1 (n3243), .A2 (n3417), .B (n1272), .Y (y1412) );
  AND3x1_ASAP7_75t_R   g3411( .A (n382), .B (y3377), .C (n724), .Y (y2612) );
  AND2x2_ASAP7_75t_R   g3412( .A (y2612), .B (x0), .Y (y1413) );
  AO21x1_ASAP7_75t_R   g3413( .A1 (n1000), .A2 (x0), .B (n1095), .Y (y1414) );
  AND3x1_ASAP7_75t_R   g3414( .A (n2542), .B (n1272), .C (n556), .Y (y1415) );
  AND3x1_ASAP7_75t_R   g3415( .A (n12), .B (n22), .C (x1), .Y (n3423) );
  INVx1_ASAP7_75t_R    g3416( .A (n3423), .Y (n3424) );
  AND2x2_ASAP7_75t_R   g3417( .A (n3380), .B (n3424), .Y (y1416) );
  NAND2x1_ASAP7_75t_R  g3418( .A (x5), .B (n415), .Y (n3426) );
  AND3x1_ASAP7_75t_R   g3419( .A (n363), .B (n22), .C (n17), .Y (n3427) );
  INVx1_ASAP7_75t_R    g3420( .A (n3427), .Y (n3428) );
  OA21x2_ASAP7_75t_R   g3421( .A1 (n2994), .A2 (n3426), .B (n3428), .Y (y1417) );
  OR3x1_ASAP7_75t_R    g3422( .A (n45), .B (x4), .C (x5), .Y (n3430) );
  AND2x2_ASAP7_75t_R   g3423( .A (n3430), .B (y3293), .Y (y1418) );
  AND2x2_ASAP7_75t_R   g3424( .A (n2688), .B (n52), .Y (y1419) );
  AO21x1_ASAP7_75t_R   g3425( .A1 (n12), .A2 (x1), .B (n518), .Y (n3433) );
  NOR2x1_ASAP7_75t_R   g3426( .A (x4), .B (n488), .Y (n3434) );
  NOR2x1_ASAP7_75t_R   g3427( .A (n3433), .B (n3434), .Y (y1420) );
  AND3x1_ASAP7_75t_R   g3428( .A (n125), .B (y2079), .C (n22), .Y (n3436) );
  NOR2x1_ASAP7_75t_R   g3429( .A (n518), .B (n3436), .Y (y1421) );
  AO21x1_ASAP7_75t_R   g3430( .A1 (n16), .A2 (n925), .B (y2826), .Y (y1422) );
  AO21x1_ASAP7_75t_R   g3431( .A1 (n12), .A2 (x3), .B (n392), .Y (n3439) );
  INVx1_ASAP7_75t_R    g3432( .A (n3439), .Y (y1423) );
  OA21x2_ASAP7_75t_R   g3433( .A1 (y3758), .A2 (n84), .B (n1620), .Y (y1424) );
  NAND2x1_ASAP7_75t_R  g3434( .A (n3160), .B (n310), .Y (y1425) );
  AND3x1_ASAP7_75t_R   g3435( .A (y2079), .B (x4), .C (x3), .Y (n3443) );
  AO21x1_ASAP7_75t_R   g3436( .A1 (n3387), .A2 (n3128), .B (n3443), .Y (y1426) );
  AO21x1_ASAP7_75t_R   g3437( .A1 (n17), .A2 (n15), .B (x4), .Y (n3445) );
  NAND2x1_ASAP7_75t_R  g3438( .A (x5), .B (n3445), .Y (n3446) );
  AND3x1_ASAP7_75t_R   g3439( .A (n22), .B (x2), .C (x3), .Y (n3447) );
  INVx1_ASAP7_75t_R    g3440( .A (n3447), .Y (n3448) );
  AND2x2_ASAP7_75t_R   g3441( .A (n3446), .B (n3448), .Y (y1427) );
  INVx1_ASAP7_75t_R    g3442( .A (n3366), .Y (n3450) );
  AO21x1_ASAP7_75t_R   g3443( .A1 (n463), .A2 (x0), .B (n3450), .Y (y1428) );
  AND2x2_ASAP7_75t_R   g3444( .A (n1755), .B (n387), .Y (y1429) );
  AND3x1_ASAP7_75t_R   g3445( .A (n63), .B (n64), .C (n1466), .Y (n3453) );
  AO21x1_ASAP7_75t_R   g3446( .A1 (n1676), .A2 (y2079), .B (n3453), .Y (y1430) );
  NAND2x1_ASAP7_75t_R  g3447( .A (n388), .B (n436), .Y (n3455) );
  AO21x1_ASAP7_75t_R   g3448( .A1 (n3455), .A2 (x0), .B (n3450), .Y (y1431) );
  AO21x1_ASAP7_75t_R   g3449( .A1 (n22), .A2 (y2079), .B (x3), .Y (n3457) );
  AO32x1_ASAP7_75t_R   g3450( .A1 (n556), .A2 (n1062), .A3 (n3457), .B1 (n15), .B2 (n455), .Y (n3458) );
  OR3x1_ASAP7_75t_R    g3451( .A (y2466), .B (n17), .C (x2), .Y (n3459) );
  AND2x2_ASAP7_75t_R   g3452( .A (n3458), .B (n3459), .Y (y1432) );
  NOR2x1_ASAP7_75t_R   g3453( .A (n58), .B (n1011), .Y (n3461) );
  NOR2x1_ASAP7_75t_R   g3454( .A (n1245), .B (n3461), .Y (n3462) );
  AND2x2_ASAP7_75t_R   g3455( .A (n3462), .B (n2596), .Y (y1433) );
  AO21x1_ASAP7_75t_R   g3456( .A1 (n1838), .A2 (n22), .B (n3023), .Y (n3464) );
  OA21x2_ASAP7_75t_R   g3457( .A1 (x2), .A2 (n407), .B (n3464), .Y (y1434) );
  AO21x1_ASAP7_75t_R   g3458( .A1 (x4), .A2 (x5), .B (n12), .Y (n3466) );
  NAND2x1_ASAP7_75t_R  g3459( .A (x1), .B (n3466), .Y (n3467) );
  AND2x2_ASAP7_75t_R   g3460( .A (n2285), .B (n3467), .Y (y1435) );
  NAND2x1_ASAP7_75t_R  g3461( .A (x4), .B (n15), .Y (n3469) );
  AND2x2_ASAP7_75t_R   g3462( .A (n360), .B (n3469), .Y (n3470) );
  AO21x1_ASAP7_75t_R   g3463( .A1 (n17), .A2 (x2), .B (n403), .Y (n3471) );
  NOR2x1_ASAP7_75t_R   g3464( .A (n3029), .B (n3471), .Y (n3472) );
  AO21x1_ASAP7_75t_R   g3465( .A1 (y2079), .A2 (n3470), .B (n3472), .Y (y1436) );
  AO21x1_ASAP7_75t_R   g3466( .A1 (n17), .A2 (x4), .B (y2079), .Y (n3474) );
  AO21x1_ASAP7_75t_R   g3467( .A1 (n189), .A2 (n22), .B (n3474), .Y (n3475) );
  INVx1_ASAP7_75t_R    g3468( .A (n3475), .Y (n3476) );
  AO21x1_ASAP7_75t_R   g3469( .A1 (n360), .A2 (n290), .B (x0), .Y (n3477) );
  NOR2x1_ASAP7_75t_R   g3470( .A (x5), .B (n3477), .Y (n3478) );
  NOR2x1_ASAP7_75t_R   g3471( .A (n3476), .B (n3478), .Y (y1437) );
  AO21x1_ASAP7_75t_R   g3472( .A1 (n12), .A2 (x5), .B (x4), .Y (n3480) );
  NAND2x1_ASAP7_75t_R  g3473( .A (n3160), .B (n3480), .Y (y1438) );
  AO21x1_ASAP7_75t_R   g3474( .A1 (n22), .A2 (x3), .B (x0), .Y (n3482) );
  AND2x2_ASAP7_75t_R   g3475( .A (n406), .B (n3482), .Y (y1439) );
  AO21x1_ASAP7_75t_R   g3476( .A1 (n3455), .A2 (x0), .B (n2001), .Y (y1440) );
  AO21x1_ASAP7_75t_R   g3477( .A1 (n16), .A2 (x5), .B (n15), .Y (n3485) );
  INVx1_ASAP7_75t_R    g3478( .A (n3485), .Y (n3486) );
  AND3x1_ASAP7_75t_R   g3479( .A (y2079), .B (x0), .C (x1), .Y (n3487) );
  AO21x1_ASAP7_75t_R   g3480( .A1 (n1242), .A2 (n271), .B (n3487), .Y (n3488) );
  AO21x1_ASAP7_75t_R   g3481( .A1 (n3486), .A2 (y195), .B (n3488), .Y (y1441) );
  AND3x1_ASAP7_75t_R   g3482( .A (n15), .B (n22), .C (x3), .Y (n3490) );
  INVx1_ASAP7_75t_R    g3483( .A (n3490), .Y (n3491) );
  AND2x2_ASAP7_75t_R   g3484( .A (n72), .B (n137), .Y (n3492) );
  INVx1_ASAP7_75t_R    g3485( .A (n3492), .Y (n3493) );
  AND2x2_ASAP7_75t_R   g3486( .A (n3493), .B (n29), .Y (n3494) );
  AO21x1_ASAP7_75t_R   g3487( .A1 (y2079), .A2 (n3491), .B (n3494), .Y (y1442) );
  AO21x1_ASAP7_75t_R   g3488( .A1 (y2079), .A2 (n436), .B (n442), .Y (n3496) );
  OR3x1_ASAP7_75t_R    g3489( .A (n544), .B (x4), .C (x0), .Y (n3497) );
  INVx1_ASAP7_75t_R    g3490( .A (n3497), .Y (n3498) );
  AO21x1_ASAP7_75t_R   g3491( .A1 (n3496), .A2 (x0), .B (n3498), .Y (y1443) );
  AO21x1_ASAP7_75t_R   g3492( .A1 (x2), .A2 (n978), .B (y890), .Y (y1444) );
  OA21x2_ASAP7_75t_R   g3493( .A1 (n518), .A2 (n3121), .B (y1903), .Y (y1446) );
  INVx1_ASAP7_75t_R    g3494( .A (n3466), .Y (n3502) );
  OA21x2_ASAP7_75t_R   g3495( .A1 (n3502), .A2 (n552), .B (n1218), .Y (y1447) );
  OR3x1_ASAP7_75t_R    g3496( .A (n143), .B (x4), .C (x5), .Y (n3504) );
  AND2x2_ASAP7_75t_R   g3497( .A (n3504), .B (y117), .Y (y1448) );
  OA21x2_ASAP7_75t_R   g3498( .A1 (n3502), .A2 (n552), .B (n1211), .Y (y1449) );
  AO21x1_ASAP7_75t_R   g3499( .A1 (n465), .A2 (x0), .B (n2001), .Y (y1450) );
  AND2x2_ASAP7_75t_R   g3500( .A (n2728), .B (n64), .Y (n3508) );
  NOR2x1_ASAP7_75t_R   g3501( .A (x3), .B (n610), .Y (n3509) );
  OA21x2_ASAP7_75t_R   g3502( .A1 (n3508), .A2 (n3509), .B (n2720), .Y (y1451) );
  AO21x1_ASAP7_75t_R   g3503( .A1 (y2079), .A2 (n401), .B (n638), .Y (n3511) );
  AO21x1_ASAP7_75t_R   g3504( .A1 (n290), .A2 (n3207), .B (x2), .Y (n3512) );
  INVx1_ASAP7_75t_R    g3505( .A (n3512), .Y (n3513) );
  AO21x1_ASAP7_75t_R   g3506( .A1 (n3511), .A2 (x2), .B (n3513), .Y (y1452) );
  AO21x1_ASAP7_75t_R   g3507( .A1 (y2079), .A2 (x0), .B (n527), .Y (n3515) );
  OA21x2_ASAP7_75t_R   g3508( .A1 (n914), .A2 (n3515), .B (n1218), .Y (y1453) );
  AO32x1_ASAP7_75t_R   g3509( .A1 (n15), .A2 (n22), .A3 (n319), .B1 (x2), .B2 (n3511), .Y (y1454) );
  AND2x2_ASAP7_75t_R   g3510( .A (y710), .B (y3293), .Y (y1455) );
  INVx1_ASAP7_75t_R    g3511( .A (n3327), .Y (n3519) );
  AO21x1_ASAP7_75t_R   g3512( .A1 (n12), .A2 (x3), .B (n22), .Y (n3520) );
  INVx1_ASAP7_75t_R    g3513( .A (n3520), .Y (n3521) );
  NOR2x1_ASAP7_75t_R   g3514( .A (n3519), .B (n3521), .Y (y1456) );
  AND3x1_ASAP7_75t_R   g3515( .A (n1062), .B (n3024), .C (y2079), .Y (n3523) );
  AO21x1_ASAP7_75t_R   g3516( .A1 (n15), .A2 (n17), .B (n22), .Y (n3524) );
  AND3x1_ASAP7_75t_R   g3517( .A (n1838), .B (n3524), .C (x5), .Y (n3525) );
  OR3x1_ASAP7_75t_R    g3518( .A (x2), .B (x3), .C (x4), .Y (n3526) );
  INVx1_ASAP7_75t_R    g3519( .A (n3526), .Y (n3527) );
  OR3x1_ASAP7_75t_R    g3520( .A (n3523), .B (n3525), .C (n3527), .Y (y1457) );
  NAND2x1_ASAP7_75t_R  g3521( .A (x1), .B (n430), .Y (n3529) );
  AND3x1_ASAP7_75t_R   g3522( .A (n3529), .B (n90), .C (y3293), .Y (y1458) );
  AO21x1_ASAP7_75t_R   g3523( .A1 (n17), .A2 (n1851), .B (n293), .Y (y1459) );
  AND3x1_ASAP7_75t_R   g3524( .A (y3758), .B (n90), .C (n219), .Y (y1460) );
  AO21x1_ASAP7_75t_R   g3525( .A1 (n15), .A2 (n988), .B (n2160), .Y (y1461) );
  AO21x1_ASAP7_75t_R   g3526( .A1 (n914), .A2 (x1), .B (y2079), .Y (y2737) );
  AND2x2_ASAP7_75t_R   g3527( .A (y2737), .B (n3366), .Y (y1462) );
  AND2x2_ASAP7_75t_R   g3528( .A (y195), .B (n482), .Y (n3536) );
  AO21x1_ASAP7_75t_R   g3529( .A1 (n312), .A2 (n315), .B (n3536), .Y (y1463) );
  OA21x2_ASAP7_75t_R   g3530( .A1 (y2147), .A2 (n1166), .B (n935), .Y (y1464) );
  INVx1_ASAP7_75t_R    g3531( .A (n2415), .Y (n3539) );
  OA211x2_ASAP7_75t_R  g3532( .A1 (n3034), .A2 (n3539), .B (n2416), .C (y9), .Y (y1465) );
  NAND2x1_ASAP7_75t_R  g3533( .A (x3), .B (n934), .Y (n3541) );
  OR3x1_ASAP7_75t_R    g3534( .A (n392), .B (n12), .C (x3), .Y (n3542) );
  AND3x1_ASAP7_75t_R   g3535( .A (n3541), .B (y1894), .C (n3542), .Y (y1466) );
  INVx1_ASAP7_75t_R    g3536( .A (n608), .Y (y1467) );
  OA21x2_ASAP7_75t_R   g3537( .A1 (n25), .A2 (n315), .B (n1247), .Y (y1468) );
  AND2x2_ASAP7_75t_R   g3538( .A (y2737), .B (n453), .Y (y1469) );
  AO21x1_ASAP7_75t_R   g3539( .A1 (y2079), .A2 (y9), .B (n1150), .Y (y1470) );
  AO21x1_ASAP7_75t_R   g3540( .A1 (n22), .A2 (x5), .B (n76), .Y (n3548) );
  AO21x1_ASAP7_75t_R   g3541( .A1 (n22), .A2 (n1572), .B (n3548), .Y (n3549) );
  OR3x1_ASAP7_75t_R    g3542( .A (n671), .B (n15), .C (x4), .Y (n3550) );
  AND3x1_ASAP7_75t_R   g3543( .A (n3549), .B (n3550), .C (n369), .Y (y1471) );
  AND2x2_ASAP7_75t_R   g3544( .A (n2952), .B (x0), .Y (n3552) );
  AO21x1_ASAP7_75t_R   g3545( .A1 (x1), .A2 (n2060), .B (n3552), .Y (y1472) );
  OA21x2_ASAP7_75t_R   g3546( .A1 (n407), .A2 (n3384), .B (y1903), .Y (y1473) );
  AO21x1_ASAP7_75t_R   g3547( .A1 (x2), .A2 (n22), .B (n3023), .Y (y1474) );
  NOR2x1_ASAP7_75t_R   g3548( .A (n15), .B (n671), .Y (n3556) );
  AO32x1_ASAP7_75t_R   g3549( .A1 (n15), .A2 (n360), .A3 (n319), .B1 (n3119), .B2 (n3556), .Y (y1475) );
  NOR2x1_ASAP7_75t_R   g3550( .A (x4), .B (n1431), .Y (n3558) );
  OR3x1_ASAP7_75t_R    g3551( .A (n3558), .B (n349), .C (n58), .Y (y1476) );
  AO21x1_ASAP7_75t_R   g3552( .A1 (n1454), .A2 (n913), .B (y247), .Y (y1477) );
  AND3x1_ASAP7_75t_R   g3553( .A (n218), .B (n388), .C (n28), .Y (n3561) );
  AO21x1_ASAP7_75t_R   g3554( .A1 (y3758), .A2 (n217), .B (n3561), .Y (y1478) );
  AO21x1_ASAP7_75t_R   g3555( .A1 (x4), .A2 (n15), .B (n319), .Y (n3563) );
  INVx1_ASAP7_75t_R    g3556( .A (n3563), .Y (n3564) );
  AO21x1_ASAP7_75t_R   g3557( .A1 (x3), .A2 (x4), .B (y2079), .Y (n3565) );
  AND3x1_ASAP7_75t_R   g3558( .A (n401), .B (n757), .C (n3565), .Y (n3566) );
  NAND2x1_ASAP7_75t_R  g3559( .A (x2), .B (n22), .Y (n3567) );
  INVx1_ASAP7_75t_R    g3560( .A (n3567), .Y (n3568) );
  OR3x1_ASAP7_75t_R    g3561( .A (n3564), .B (n3566), .C (n3568), .Y (y1479) );
  AO21x1_ASAP7_75t_R   g3562( .A1 (n16), .A2 (x0), .B (n999), .Y (n3570) );
  NAND2x1_ASAP7_75t_R  g3563( .A (x5), .B (n1150), .Y (n3571) );
  INVx1_ASAP7_75t_R    g3564( .A (n3571), .Y (n3572) );
  AO21x1_ASAP7_75t_R   g3565( .A1 (y2079), .A2 (n3570), .B (n3572), .Y (y1480) );
  INVx1_ASAP7_75t_R    g3566( .A (n415), .Y (n3574) );
  OR3x1_ASAP7_75t_R    g3567( .A (n3574), .B (n3521), .C (y2079), .Y (y1481) );
  NAND2x1_ASAP7_75t_R  g3568( .A (n1242), .B (n436), .Y (n3576) );
  AO21x1_ASAP7_75t_R   g3569( .A1 (x0), .A2 (x5), .B (x4), .Y (n3577) );
  AND2x2_ASAP7_75t_R   g3570( .A (n3576), .B (n3577), .Y (y1482) );
  AO21x1_ASAP7_75t_R   g3571( .A1 (n12), .A2 (y2079), .B (n17), .Y (n3579) );
  INVx1_ASAP7_75t_R    g3572( .A (n3579), .Y (n3580) );
  NAND2x1_ASAP7_75t_R  g3573( .A (x3), .B (n614), .Y (n3581) );
  OA21x2_ASAP7_75t_R   g3574( .A1 (n3580), .A2 (n22), .B (n3581), .Y (y1483) );
  AO21x1_ASAP7_75t_R   g3575( .A1 (y2079), .A2 (n3471), .B (n3472), .Y (y1484) );
  AO21x1_ASAP7_75t_R   g3576( .A1 (n15), .A2 (x4), .B (x5), .Y (n3584) );
  INVx1_ASAP7_75t_R    g3577( .A (n3584), .Y (n3585) );
  AO21x1_ASAP7_75t_R   g3578( .A1 (n1062), .A2 (x4), .B (n2999), .Y (n3586) );
  AO32x1_ASAP7_75t_R   g3579( .A1 (n672), .A2 (n3000), .A3 (n3524), .B1 (n3585), .B2 (n3586), .Y (y1485) );
  AO21x1_ASAP7_75t_R   g3580( .A1 (x2), .A2 (x3), .B (y2079), .Y (n3588) );
  NAND2x1_ASAP7_75t_R  g3581( .A (x4), .B (n3588), .Y (n3589) );
  AO21x1_ASAP7_75t_R   g3582( .A1 (n3588), .A2 (x4), .B (n29), .Y (n3590) );
  AO32x1_ASAP7_75t_R   g3583( .A1 (n28), .A2 (n3589), .A3 (n217), .B1 (n218), .B2 (n3590), .Y (y1486) );
  AO21x1_ASAP7_75t_R   g3584( .A1 (y2079), .A2 (n1062), .B (n2989), .Y (n3592) );
  AO21x1_ASAP7_75t_R   g3585( .A1 (n45), .A2 (n455), .B (n3592), .Y (y1487) );
  AND3x1_ASAP7_75t_R   g3586( .A (n221), .B (n137), .C (n72), .Y (n3594) );
  AO21x1_ASAP7_75t_R   g3587( .A1 (n218), .A2 (y435), .B (n3594), .Y (n3595) );
  INVx1_ASAP7_75t_R    g3588( .A (n3595), .Y (y1488) );
  AO21x1_ASAP7_75t_R   g3589( .A1 (n22), .A2 (n3191), .B (n3107), .Y (y1489) );
  AND3x1_ASAP7_75t_R   g3590( .A (x3), .B (x5), .C (x4), .Y (n3598) );
  AO21x1_ASAP7_75t_R   g3591( .A1 (n1838), .A2 (n418), .B (n3598), .Y (n3599) );
  NAND2x1_ASAP7_75t_R  g3592( .A (n295), .B (n391), .Y (n3600) );
  AND2x2_ASAP7_75t_R   g3593( .A (n3600), .B (x2), .Y (n3601) );
  AO21x1_ASAP7_75t_R   g3594( .A1 (n15), .A2 (n3599), .B (n3601), .Y (y1490) );
  NOR2x1_ASAP7_75t_R   g3595( .A (n16), .B (n537), .Y (n3603) );
  AO21x1_ASAP7_75t_R   g3596( .A1 (n299), .A2 (n310), .B (n16), .Y (n3604) );
  INVx1_ASAP7_75t_R    g3597( .A (n3604), .Y (n3605) );
  NAND2x1_ASAP7_75t_R  g3598( .A (y2079), .B (n3605), .Y (n3606) );
  OA211x2_ASAP7_75t_R  g3599( .A1 (n3417), .A2 (n3603), .B (n3606), .C (y3852), .Y (y1491) );
  NOR2x1_ASAP7_75t_R   g3600( .A (x5), .B (n2980), .Y (n3608) );
  INVx1_ASAP7_75t_R    g3601( .A (n3608), .Y (n3609) );
  AND2x2_ASAP7_75t_R   g3602( .A (n3609), .B (n3030), .Y (y1492) );
  AND3x1_ASAP7_75t_R   g3603( .A (y2079), .B (x3), .C (x2), .Y (n3611) );
  INVx1_ASAP7_75t_R    g3604( .A (n3611), .Y (n3612) );
  AO21x1_ASAP7_75t_R   g3605( .A1 (n3612), .A2 (n1062), .B (n22), .Y (n3613) );
  OAI21x1_ASAP7_75t_R  g3606( .A1 (n3294), .A2 (n3024), .B (n3613), .Y (y1493) );
  AO21x1_ASAP7_75t_R   g3607( .A1 (n71), .A2 (n69), .B (n103), .Y (y1494) );
  AO21x1_ASAP7_75t_R   g3608( .A1 (n16), .A2 (n572), .B (n1140), .Y (y1495) );
  AND3x1_ASAP7_75t_R   g3609( .A (n15), .B (x4), .C (x5), .Y (n3617) );
  AO21x1_ASAP7_75t_R   g3610( .A1 (n15), .A2 (n22), .B (n17), .Y (n3618) );
  OA22x2_ASAP7_75t_R   g3611( .A1 (n3617), .A2 (n3181), .B1 (n1269), .B2 (n3618), .Y (y1496) );
  AO21x1_ASAP7_75t_R   g3612( .A1 (n22), .A2 (x3), .B (n12), .Y (n3620) );
  AND3x1_ASAP7_75t_R   g3613( .A (n84), .B (n3620), .C (y2079), .Y (n3621) );
  INVx1_ASAP7_75t_R    g3614( .A (n3621), .Y (n3622) );
  AND2x2_ASAP7_75t_R   g3615( .A (n3622), .B (y1343), .Y (y1497) );
  AND3x1_ASAP7_75t_R   g3616( .A (n856), .B (n22), .C (n17), .Y (n3624) );
  INVx1_ASAP7_75t_R    g3617( .A (n3624), .Y (n3625) );
  AO21x1_ASAP7_75t_R   g3618( .A1 (n15), .A2 (y2079), .B (n22), .Y (n3626) );
  AND3x1_ASAP7_75t_R   g3619( .A (n3625), .B (n3626), .C (n369), .Y (y1498) );
  NOR2x1_ASAP7_75t_R   g3620( .A (n3027), .B (n319), .Y (n3628) );
  AO21x1_ASAP7_75t_R   g3621( .A1 (x2), .A2 (x4), .B (x3), .Y (n3629) );
  AO21x1_ASAP7_75t_R   g3622( .A1 (y2079), .A2 (x2), .B (n2999), .Y (n3630) );
  AO32x1_ASAP7_75t_R   g3623( .A1 (n3000), .A2 (n3628), .A3 (n740), .B1 (n3629), .B2 (n3630), .Y (y1499) );
  AND2x2_ASAP7_75t_R   g3624( .A (n1969), .B (x0), .Y (n3632) );
  AO21x1_ASAP7_75t_R   g3625( .A1 (n2017), .A2 (n16), .B (n3632), .Y (y1500) );
  AND3x1_ASAP7_75t_R   g3626( .A (n84), .B (n3128), .C (x5), .Y (n3634) );
  AO21x1_ASAP7_75t_R   g3627( .A1 (x3), .A2 (n529), .B (n3634), .Y (y1501) );
  AO21x1_ASAP7_75t_R   g3628( .A1 (y2079), .A2 (x3), .B (x2), .Y (n3636) );
  INVx1_ASAP7_75t_R    g3629( .A (n3469), .Y (n3637) );
  AND2x2_ASAP7_75t_R   g3630( .A (n316), .B (n319), .Y (n3638) );
  AO221x2_ASAP7_75t_R  g3631( .A1 (n3284), .A2 (n3636), .B1 (n3637), .B2 (n3638), .C (n1269), .Y (y1502) );
  AO21x1_ASAP7_75t_R   g3632( .A1 (n583), .A2 (n22), .B (n3360), .Y (n3640) );
  INVx1_ASAP7_75t_R    g3633( .A (n3640), .Y (n3641) );
  AO21x1_ASAP7_75t_R   g3634( .A1 (n17), .A2 (y1467), .B (n3641), .Y (n3642) );
  NAND2x1_ASAP7_75t_R  g3635( .A (n622), .B (n3642), .Y (y1503) );
  OR3x1_ASAP7_75t_R    g3636( .A (n529), .B (n3568), .C (n45), .Y (y1504) );
  AO21x1_ASAP7_75t_R   g3637( .A1 (y2079), .A2 (x0), .B (n17), .Y (n3645) );
  INVx1_ASAP7_75t_R    g3638( .A (n3645), .Y (n3646) );
  NAND2x1_ASAP7_75t_R  g3639( .A (x4), .B (n3646), .Y (n3647) );
  OR3x1_ASAP7_75t_R    g3640( .A (n518), .B (n12), .C (x3), .Y (n3648) );
  AO21x1_ASAP7_75t_R   g3641( .A1 (n3648), .A2 (n652), .B (y2079), .Y (n3649) );
  AND2x2_ASAP7_75t_R   g3642( .A (n3647), .B (n3649), .Y (y1505) );
  OR3x1_ASAP7_75t_R    g3643( .A (n982), .B (n914), .C (n529), .Y (y1506) );
  AND3x1_ASAP7_75t_R   g3644( .A (n12), .B (n17), .C (x2), .Y (n3652) );
  OR3x1_ASAP7_75t_R    g3645( .A (n2588), .B (n3652), .C (n73), .Y (y1507) );
  AND2x2_ASAP7_75t_R   g3646( .A (n3606), .B (y2737), .Y (y1508) );
  OR3x1_ASAP7_75t_R    g3647( .A (n163), .B (n164), .C (n3207), .Y (n3655) );
  AND2x2_ASAP7_75t_R   g3648( .A (n3655), .B (n556), .Y (y1509) );
  AND2x2_ASAP7_75t_R   g3649( .A (n3284), .B (x2), .Y (n3657) );
  AO21x1_ASAP7_75t_R   g3650( .A1 (n3183), .A2 (x3), .B (n3657), .Y (y1510) );
  AND3x1_ASAP7_75t_R   g3651( .A (n22), .B (n17), .C (x2), .Y (n3659) );
  INVx1_ASAP7_75t_R    g3652( .A (n3659), .Y (n3660) );
  NAND2x1_ASAP7_75t_R  g3653( .A (y2079), .B (n2980), .Y (n3661) );
  INVx1_ASAP7_75t_R    g3654( .A (n3661), .Y (n3662) );
  AO21x1_ASAP7_75t_R   g3655( .A1 (n3660), .A2 (n288), .B (n3662), .Y (y1511) );
  AO21x1_ASAP7_75t_R   g3656( .A1 (n437), .A2 (y3852), .B (n990), .Y (y1512) );
  AND2x2_ASAP7_75t_R   g3657( .A (n1188), .B (n463), .Y (y1513) );
  AO21x1_ASAP7_75t_R   g3658( .A1 (x5), .A2 (n12), .B (n436), .Y (n3666) );
  INVx1_ASAP7_75t_R    g3659( .A (n3666), .Y (n3667) );
  AO21x1_ASAP7_75t_R   g3660( .A1 (y2079), .A2 (n1077), .B (n3667), .Y (y1514) );
  AND2x2_ASAP7_75t_R   g3661( .A (n463), .B (x0), .Y (y1515) );
  AO21x1_ASAP7_75t_R   g3662( .A1 (n189), .A2 (n660), .B (n2184), .Y (y1516) );
  AND2x2_ASAP7_75t_R   g3663( .A (y563), .B (n546), .Y (y1517) );
  AO21x1_ASAP7_75t_R   g3664( .A1 (n3455), .A2 (x0), .B (n1757), .Y (y1518) );
  AND2x2_ASAP7_75t_R   g3665( .A (n1201), .B (n1932), .Y (y1519) );
  AND3x1_ASAP7_75t_R   g3666( .A (n377), .B (n451), .C (y1281), .Y (y1520) );
  AND2x2_ASAP7_75t_R   g3667( .A (n1047), .B (n463), .Y (y3447) );
  AND2x2_ASAP7_75t_R   g3668( .A (n1863), .B (y3447), .Y (y1521) );
  AO21x1_ASAP7_75t_R   g3669( .A1 (n17), .A2 (n15), .B (n518), .Y (n3677) );
  OR3x1_ASAP7_75t_R    g3670( .A (n529), .B (n29), .C (n76), .Y (n3678) );
  NAND2x1_ASAP7_75t_R  g3671( .A (n3677), .B (n3678), .Y (y1522) );
  AND3x1_ASAP7_75t_R   g3672( .A (n1863), .B (n1175), .C (y2737), .Y (y1523) );
  OR3x1_ASAP7_75t_R    g3673( .A (y863), .B (x4), .C (x5), .Y (n3681) );
  AND2x2_ASAP7_75t_R   g3674( .A (n3681), .B (y1242), .Y (y1524) );
  OA21x2_ASAP7_75t_R   g3675( .A1 (n241), .A2 (x1), .B (y2079), .Y (n3683) );
  AO21x1_ASAP7_75t_R   g3676( .A1 (n824), .A2 (x0), .B (n3683), .Y (y1525) );
  AO21x1_ASAP7_75t_R   g3677( .A1 (n22), .A2 (x2), .B (n17), .Y (n3685) );
  AND3x1_ASAP7_75t_R   g3678( .A (n3660), .B (n3630), .C (n3685), .Y (y1526) );
  AO21x1_ASAP7_75t_R   g3679( .A1 (n22), .A2 (x5), .B (n990), .Y (n3687) );
  INVx1_ASAP7_75t_R    g3680( .A (n3687), .Y (n3688) );
  OR3x1_ASAP7_75t_R    g3681( .A (n529), .B (n29), .C (n2718), .Y (y3352) );
  OA21x2_ASAP7_75t_R   g3682( .A1 (n3688), .A2 (x3), .B (y3352), .Y (y1527) );
  OA21x2_ASAP7_75t_R   g3683( .A1 (n3667), .A2 (y2196), .B (n451), .Y (y1528) );
  AND2x2_ASAP7_75t_R   g3684( .A (n436), .B (n299), .Y (n3692) );
  AO21x1_ASAP7_75t_R   g3685( .A1 (y2079), .A2 (n3692), .B (n3572), .Y (y1529) );
  AND3x1_ASAP7_75t_R   g3686( .A (n22), .B (y2079), .C (x2), .Y (n3694) );
  NOR2x1_ASAP7_75t_R   g3687( .A (n3694), .B (n678), .Y (y1530) );
  AO21x1_ASAP7_75t_R   g3688( .A1 (n12), .A2 (n16), .B (n544), .Y (n3696) );
  AO21x1_ASAP7_75t_R   g3689( .A1 (n22), .A2 (n3696), .B (n493), .Y (y1531) );
  AND3x1_ASAP7_75t_R   g3690( .A (n546), .B (n463), .C (x0), .Y (y1532) );
  AO21x1_ASAP7_75t_R   g3691( .A1 (n144), .A2 (n1646), .B (n2156), .Y (y1533) );
  AND3x1_ASAP7_75t_R   g3692( .A (n12), .B (x4), .C (x1), .Y (n3700) );
  NOR2x1_ASAP7_75t_R   g3693( .A (x5), .B (n3700), .Y (n3701) );
  AO21x1_ASAP7_75t_R   g3694( .A1 (x5), .A2 (n16), .B (n310), .Y (n3702) );
  INVx1_ASAP7_75t_R    g3695( .A (n3702), .Y (n3703) );
  AO21x1_ASAP7_75t_R   g3696( .A1 (n719), .A2 (n3701), .B (n3703), .Y (y1534) );
  INVx1_ASAP7_75t_R    g3697( .A (n2989), .Y (n3705) );
  AO21x1_ASAP7_75t_R   g3698( .A1 (n3705), .A2 (n3469), .B (x5), .Y (n3706) );
  OR3x1_ASAP7_75t_R    g3699( .A (n2989), .B (y2079), .C (n45), .Y (y3171) );
  AND2x2_ASAP7_75t_R   g3700( .A (n3706), .B (y3171), .Y (y1535) );
  AND3x1_ASAP7_75t_R   g3701( .A (n90), .B (n219), .C (n463), .Y (y1536) );
  AND3x1_ASAP7_75t_R   g3702( .A (n382), .B (y3377), .C (x2), .Y (n3710) );
  NOR2x1_ASAP7_75t_R   g3703( .A (n3218), .B (n3710), .Y (y1537) );
  OR3x1_ASAP7_75t_R    g3704( .A (n1205), .B (y2079), .C (n537), .Y (n3712) );
  OR3x1_ASAP7_75t_R    g3705( .A (n1208), .B (n596), .C (x5), .Y (n3713) );
  AND2x2_ASAP7_75t_R   g3706( .A (n3712), .B (n3713), .Y (y1538) );
  AO21x1_ASAP7_75t_R   g3707( .A1 (x1), .A2 (x0), .B (n950), .Y (n3715) );
  AND2x2_ASAP7_75t_R   g3708( .A (n3715), .B (n556), .Y (y1539) );
  NOR2x1_ASAP7_75t_R   g3709( .A (n518), .B (n2989), .Y (y1540) );
  OR3x1_ASAP7_75t_R    g3710( .A (n756), .B (n22), .C (n17), .Y (n3718) );
  INVx1_ASAP7_75t_R    g3711( .A (n3718), .Y (n3719) );
  AO21x1_ASAP7_75t_R   g3712( .A1 (n97), .A2 (n3284), .B (n3719), .Y (y1541) );
  AO21x1_ASAP7_75t_R   g3713( .A1 (n276), .A2 (x1), .B (n17), .Y (n3721) );
  OA21x2_ASAP7_75t_R   g3714( .A1 (n43), .A2 (n137), .B (n3721), .Y (y1542) );
  AND3x1_ASAP7_75t_R   g3715( .A (n1676), .B (y2079), .C (x0), .Y (n3723) );
  INVx1_ASAP7_75t_R    g3716( .A (n3723), .Y (n3724) );
  AND2x2_ASAP7_75t_R   g3717( .A (n3724), .B (y238), .Y (y1543) );
  AND3x1_ASAP7_75t_R   g3718( .A (n189), .B (n310), .C (y2079), .Y (n3726) );
  AO21x1_ASAP7_75t_R   g3719( .A1 (n22), .A2 (n3191), .B (n3726), .Y (y1544) );
  AND3x1_ASAP7_75t_R   g3720( .A (n3195), .B (n546), .C (n387), .Y (y1545) );
  OA21x2_ASAP7_75t_R   g3721( .A1 (y3758), .A2 (n1208), .B (y3852), .Y (y1546) );
  NOR2x1_ASAP7_75t_R   g3722( .A (n450), .B (n1927), .Y (y1891) );
  AND3x1_ASAP7_75t_R   g3723( .A (y1891), .B (n90), .C (n219), .Y (y1547) );
  AND3x1_ASAP7_75t_R   g3724( .A (n22), .B (x0), .C (x1), .Y (n3732) );
  AO21x1_ASAP7_75t_R   g3725( .A1 (n1240), .A2 (y2079), .B (n3732), .Y (y1548) );
  AO21x1_ASAP7_75t_R   g3726( .A1 (n22), .A2 (n77), .B (n3132), .Y (y2016) );
  AND2x2_ASAP7_75t_R   g3727( .A (y2016), .B (n1572), .Y (y1549) );
  AO21x1_ASAP7_75t_R   g3728( .A1 (n84), .A2 (n125), .B (x4), .Y (n3736) );
  AND3x1_ASAP7_75t_R   g3729( .A (y1903), .B (n3736), .C (n672), .Y (y1550) );
  OR3x1_ASAP7_75t_R    g3730( .A (y863), .B (x5), .C (x4), .Y (n3738) );
  NAND2x1_ASAP7_75t_R  g3731( .A (n1744), .B (n3738), .Y (n3739) );
  OA21x2_ASAP7_75t_R   g3732( .A1 (n914), .A2 (n495), .B (n3739), .Y (y1551) );
  AO21x1_ASAP7_75t_R   g3733( .A1 (n16), .A2 (x0), .B (n392), .Y (n3741) );
  INVx1_ASAP7_75t_R    g3734( .A (n3741), .Y (n3742) );
  AO21x1_ASAP7_75t_R   g3735( .A1 (n3742), .A2 (n469), .B (n1399), .Y (y1552) );
  OR3x1_ASAP7_75t_R    g3736( .A (n392), .B (n16), .C (n12), .Y (n3744) );
  INVx1_ASAP7_75t_R    g3737( .A (n3744), .Y (y3160) );
  OA21x2_ASAP7_75t_R   g3738( .A1 (y3160), .A2 (n418), .B (n469), .Y (y1554) );
  NOR2x1_ASAP7_75t_R   g3739( .A (n1980), .B (n43), .Y (n3747) );
  INVx1_ASAP7_75t_R    g3740( .A (y250), .Y (n3748) );
  NOR2x1_ASAP7_75t_R   g3741( .A (n3747), .B (n3748), .Y (y1555) );
  AND2x2_ASAP7_75t_R   g3742( .A (n1062), .B (n3567), .Y (n3750) );
  NOR2x1_ASAP7_75t_R   g3743( .A (y2079), .B (n3750), .Y (n3751) );
  AO21x1_ASAP7_75t_R   g3744( .A1 (y2079), .A2 (n3750), .B (n3751), .Y (y1556) );
  OR3x1_ASAP7_75t_R    g3745( .A (n1770), .B (n1817), .C (n143), .Y (y1557) );
  OR3x1_ASAP7_75t_R    g3746( .A (n529), .B (n29), .C (n43), .Y (n3754) );
  AO21x1_ASAP7_75t_R   g3747( .A1 (n22), .A2 (y2079), .B (n143), .Y (n3755) );
  AND2x2_ASAP7_75t_R   g3748( .A (n3754), .B (n3755), .Y (y1558) );
  AND3x1_ASAP7_75t_R   g3749( .A (n1196), .B (n219), .C (n419), .Y (y1559) );
  AO21x1_ASAP7_75t_R   g3750( .A1 (n1851), .A2 (n628), .B (n3257), .Y (y1560) );
  AND2x2_ASAP7_75t_R   g3751( .A (n806), .B (n2276), .Y (y1561) );
  AO21x1_ASAP7_75t_R   g3752( .A1 (x3), .A2 (n22), .B (n3474), .Y (y1693) );
  INVx1_ASAP7_75t_R    g3753( .A (y1693), .Y (n3761) );
  AO21x1_ASAP7_75t_R   g3754( .A1 (n17), .A2 (n22), .B (x2), .Y (n3762) );
  INVx1_ASAP7_75t_R    g3755( .A (n3762), .Y (n3763) );
  AOI22x1_ASAP7_75t_R  g3756( .A1 (n3761), .A2 (n3762), .B1 (n3763), .B2 (y1693), .Y (y1562) );
  AO21x1_ASAP7_75t_R   g3757( .A1 (n466), .A2 (n219), .B (n1817), .Y (y1563) );
  AO21x1_ASAP7_75t_R   g3758( .A1 (n388), .A2 (n28), .B (n12), .Y (n3766) );
  NOR2x1_ASAP7_75t_R   g3759( .A (n16), .B (n3766), .Y (y1564) );
  AO21x1_ASAP7_75t_R   g3760( .A1 (n2718), .A2 (n22), .B (y2079), .Y (y3198) );
  AND2x2_ASAP7_75t_R   g3761( .A (y3198), .B (n660), .Y (y1876) );
  AOI21x1_ASAP7_75t_R  g3762( .A1 (n3072), .A2 (n3519), .B (y1876), .Y (y1565) );
  AO21x1_ASAP7_75t_R   g3763( .A1 (n3124), .A2 (n1838), .B (n3099), .Y (y1566) );
  AND2x2_ASAP7_75t_R   g3764( .A (n1891), .B (n387), .Y (y1567) );
  AND2x2_ASAP7_75t_R   g3765( .A (n1974), .B (n1272), .Y (y1568) );
  NOR2x1_ASAP7_75t_R   g3766( .A (x5), .B (n2999), .Y (n3774) );
  AO21x1_ASAP7_75t_R   g3767( .A1 (n29), .A2 (n1838), .B (n3774), .Y (y1569) );
  AO21x1_ASAP7_75t_R   g3768( .A1 (n17), .A2 (y2079), .B (x4), .Y (n3776) );
  INVx1_ASAP7_75t_R    g3769( .A (n3776), .Y (n3777) );
  NAND2x1_ASAP7_75t_R  g3770( .A (x5), .B (n3620), .Y (n3778) );
  OA21x2_ASAP7_75t_R   g3771( .A1 (n3777), .A2 (n12), .B (n3778), .Y (y1570) );
  AO21x1_ASAP7_75t_R   g3772( .A1 (x5), .A2 (x4), .B (n15), .Y (n3780) );
  INVx1_ASAP7_75t_R    g3773( .A (n3780), .Y (n3781) );
  AO21x1_ASAP7_75t_R   g3774( .A1 (x5), .A2 (n3263), .B (n3781), .Y (y1571) );
  AO21x1_ASAP7_75t_R   g3775( .A1 (n645), .A2 (n3327), .B (n378), .Y (y1572) );
  AND3x1_ASAP7_75t_R   g3776( .A (n90), .B (n219), .C (x4), .Y (n3784) );
  NAND2x1_ASAP7_75t_R  g3777( .A (x5), .B (n3732), .Y (n3785) );
  INVx1_ASAP7_75t_R    g3778( .A (n3785), .Y (n3786) );
  AO21x1_ASAP7_75t_R   g3779( .A1 (y2079), .A2 (n3784), .B (n3786), .Y (y1573) );
  AO21x1_ASAP7_75t_R   g3780( .A1 (n2298), .A2 (n1490), .B (y2079), .Y (y1574) );
  NAND2x1_ASAP7_75t_R  g3781( .A (n22), .B (n2971), .Y (n3789) );
  OR3x1_ASAP7_75t_R    g3782( .A (n3447), .B (y2079), .C (n81), .Y (n3790) );
  OA21x2_ASAP7_75t_R   g3783( .A1 (n218), .A2 (n3789), .B (n3790), .Y (y1575) );
  AO21x1_ASAP7_75t_R   g3784( .A1 (n12), .A2 (n17), .B (n403), .Y (n3792) );
  OA21x2_ASAP7_75t_R   g3785( .A1 (n3792), .A2 (n58), .B (n556), .Y (y1576) );
  AO21x1_ASAP7_75t_R   g3786( .A1 (n17), .A2 (n15), .B (x5), .Y (n3794) );
  AO21x1_ASAP7_75t_R   g3787( .A1 (n3794), .A2 (n3316), .B (n529), .Y (y1577) );
  AND3x1_ASAP7_75t_R   g3788( .A (y2466), .B (n17), .C (x0), .Y (n3796) );
  INVx1_ASAP7_75t_R    g3789( .A (n3796), .Y (n3797) );
  AND3x1_ASAP7_75t_R   g3790( .A (n3797), .B (n718), .C (n369), .Y (y1578) );
  AO21x1_ASAP7_75t_R   g3791( .A1 (n2577), .A2 (y9), .B (n15), .Y (n3799) );
  AO21x1_ASAP7_75t_R   g3792( .A1 (x0), .A2 (x1), .B (n17), .Y (n3800) );
  OA211x2_ASAP7_75t_R  g3793( .A1 (n1635), .A2 (n2576), .B (n3799), .C (n3800), .Y (y1579) );
  INVx1_ASAP7_75t_R    g3794( .A (n2828), .Y (n3802) );
  OA21x2_ASAP7_75t_R   g3795( .A1 (n3802), .A2 (x4), .B (n556), .Y (y1580) );
  AO21x1_ASAP7_75t_R   g3796( .A1 (n17), .A2 (n15), .B (n22), .Y (n3804) );
  NAND2x1_ASAP7_75t_R  g3797( .A (y2079), .B (n3804), .Y (n3805) );
  INVx1_ASAP7_75t_R    g3798( .A (n3805), .Y (y1581) );
  AO21x1_ASAP7_75t_R   g3799( .A1 (x0), .A2 (x2), .B (x5), .Y (n3807) );
  INVx1_ASAP7_75t_R    g3800( .A (n3807), .Y (n3808) );
  AO21x1_ASAP7_75t_R   g3801( .A1 (n63), .A2 (n3808), .B (n530), .Y (y1582) );
  AO21x1_ASAP7_75t_R   g3802( .A1 (n290), .A2 (n360), .B (x2), .Y (n3810) );
  INVx1_ASAP7_75t_R    g3803( .A (n3810), .Y (n3811) );
  AOI22x1_ASAP7_75t_R  g3804( .A1 (n3811), .A2 (n366), .B1 (n3301), .B2 (n3810), .Y (y1583) );
  OA21x2_ASAP7_75t_R   g3805( .A1 (n529), .A2 (n661), .B (n642), .Y (y1584) );
  OR3x1_ASAP7_75t_R    g3806( .A (n987), .B (n1004), .C (n143), .Y (y1585) );
  AND3x1_ASAP7_75t_R   g3807( .A (n1971), .B (n219), .C (n455), .Y (y1586) );
  AO21x1_ASAP7_75t_R   g3808( .A1 (y2079), .A2 (n1707), .B (n3732), .Y (y1587) );
  AO21x1_ASAP7_75t_R   g3809( .A1 (y2079), .A2 (x2), .B (x4), .Y (n3817) );
  INVx1_ASAP7_75t_R    g3810( .A (n3817), .Y (n3818) );
  AND3x1_ASAP7_75t_R   g3811( .A (y2079), .B (x4), .C (x2), .Y (n3819) );
  OA21x2_ASAP7_75t_R   g3812( .A1 (n3818), .A2 (n3819), .B (n17), .Y (n3820) );
  AO21x1_ASAP7_75t_R   g3813( .A1 (n3028), .A2 (n628), .B (n3820), .Y (y1588) );
  NAND2x1_ASAP7_75t_R  g3814( .A (n3282), .B (n3794), .Y (y1589) );
  AO21x1_ASAP7_75t_R   g3815( .A1 (y2079), .A2 (n22), .B (x2), .Y (n3823) );
  NAND2x1_ASAP7_75t_R  g3816( .A (n17), .B (n3823), .Y (n3824) );
  OR3x1_ASAP7_75t_R    g3817( .A (n418), .B (n17), .C (x2), .Y (n3825) );
  AND3x1_ASAP7_75t_R   g3818( .A (n3824), .B (n3825), .C (n3780), .Y (n3826) );
  INVx1_ASAP7_75t_R    g3819( .A (n3826), .Y (y1590) );
  AO21x1_ASAP7_75t_R   g3820( .A1 (n15), .A2 (x5), .B (n17), .Y (n3828) );
  NAND2x1_ASAP7_75t_R  g3821( .A (y2079), .B (n3143), .Y (n3829) );
  INVx1_ASAP7_75t_R    g3822( .A (n3829), .Y (n3830) );
  AO21x1_ASAP7_75t_R   g3823( .A1 (n22), .A2 (n3828), .B (n3830), .Y (y1591) );
  OR3x1_ASAP7_75t_R    g3824( .A (x3), .B (x5), .C (x4), .Y (n3832) );
  AND3x1_ASAP7_75t_R   g3825( .A (n3014), .B (n3832), .C (n15), .Y (n3833) );
  INVx1_ASAP7_75t_R    g3826( .A (n3833), .Y (n3834) );
  OR3x1_ASAP7_75t_R    g3827( .A (n418), .B (n17), .C (n15), .Y (n3835) );
  AND3x1_ASAP7_75t_R   g3828( .A (n3834), .B (n3835), .C (y3293), .Y (y1592) );
  NAND2x1_ASAP7_75t_R  g3829( .A (x2), .B (n3014), .Y (n3837) );
  AOI21x1_ASAP7_75t_R  g3830( .A1 (n3825), .A2 (n3837), .B (n392), .Y (y1593) );
  OA21x2_ASAP7_75t_R   g3831( .A1 (y1467), .A2 (x1), .B (n1040), .Y (y1594) );
  INVx1_ASAP7_75t_R    g3832( .A (n1517), .Y (n3840) );
  AO21x1_ASAP7_75t_R   g3833( .A1 (x2), .A2 (n12), .B (n626), .Y (n3841) );
  INVx1_ASAP7_75t_R    g3834( .A (n3841), .Y (n3842) );
  NAND2x1_ASAP7_75t_R  g3835( .A (n2415), .B (n3840), .Y (n3843) );
  AO32x1_ASAP7_75t_R   g3836( .A1 (n2415), .A2 (n3840), .A3 (n3841), .B1 (n3842), .B2 (n3843), .Y (y1595) );
  AO21x1_ASAP7_75t_R   g3837( .A1 (y2079), .A2 (x2), .B (n337), .Y (n3845) );
  AO21x1_ASAP7_75t_R   g3838( .A1 (n1646), .A2 (n660), .B (n3845), .Y (y3085) );
  AND3x1_ASAP7_75t_R   g3839( .A (n337), .B (n15), .C (x5), .Y (n3847) );
  INVx1_ASAP7_75t_R    g3840( .A (n3847), .Y (n3848) );
  AND2x2_ASAP7_75t_R   g3841( .A (y3085), .B (n3848), .Y (y1596) );
  OR3x1_ASAP7_75t_R    g3842( .A (y2466), .B (n15), .C (x3), .Y (n3850) );
  OA21x2_ASAP7_75t_R   g3843( .A1 (n3298), .A2 (n1277), .B (n3850), .Y (y1597) );
  NAND2x1_ASAP7_75t_R  g3844( .A (n12), .B (n457), .Y (n3852) );
  AND2x2_ASAP7_75t_R   g3845( .A (n3852), .B (n1196), .Y (y1598) );
  NOR2x1_ASAP7_75t_R   g3846( .A (n15), .B (n145), .Y (n3854) );
  NOR2x1_ASAP7_75t_R   g3847( .A (n1549), .B (n3854), .Y (n3855) );
  AO22x1_ASAP7_75t_R   g3848( .A1 (n3855), .A2 (n1296), .B1 (n2415), .B2 (n3034), .Y (y1599) );
  AO21x1_ASAP7_75t_R   g3849( .A1 (n22), .A2 (x3), .B (x2), .Y (n3857) );
  AND2x2_ASAP7_75t_R   g3850( .A (n3209), .B (n3857), .Y (y1600) );
  INVx1_ASAP7_75t_R    g3851( .A (n2971), .Y (n3859) );
  AO21x1_ASAP7_75t_R   g3852( .A1 (x4), .A2 (x5), .B (n76), .Y (n3860) );
  OA21x2_ASAP7_75t_R   g3853( .A1 (n3859), .A2 (n3860), .B (y1267), .Y (y1601) );
  INVx1_ASAP7_75t_R    g3854( .A (n703), .Y (n3862) );
  AO21x1_ASAP7_75t_R   g3855( .A1 (n15), .A2 (n16), .B (n145), .Y (n3863) );
  AO21x1_ASAP7_75t_R   g3856( .A1 (n1296), .A2 (x2), .B (n2904), .Y (n3864) );
  OA21x2_ASAP7_75t_R   g3857( .A1 (n3862), .A2 (n3863), .B (n3864), .Y (y1602) );
  AO21x1_ASAP7_75t_R   g3858( .A1 (n15), .A2 (n17), .B (x5), .Y (n3866) );
  NOR2x1_ASAP7_75t_R   g3859( .A (n45), .B (n388), .Y (n3867) );
  AO21x1_ASAP7_75t_R   g3860( .A1 (n3866), .A2 (n3025), .B (n3867), .Y (y1603) );
  AO21x1_ASAP7_75t_R   g3861( .A1 (n913), .A2 (n2163), .B (n1778), .Y (y1604) );
  AO21x1_ASAP7_75t_R   g3862( .A1 (n3387), .A2 (n3128), .B (y2079), .Y (y2135) );
  AO21x1_ASAP7_75t_R   g3863( .A1 (n360), .A2 (n290), .B (n352), .Y (n3871) );
  AND2x2_ASAP7_75t_R   g3864( .A (y2135), .B (n3871), .Y (y1605) );
  AO21x1_ASAP7_75t_R   g3865( .A1 (n968), .A2 (n970), .B (n1805), .Y (y1606) );
  NAND2x1_ASAP7_75t_R  g3866( .A (n17), .B (n430), .Y (n3874) );
  OA21x2_ASAP7_75t_R   g3867( .A1 (n3874), .A2 (n3149), .B (n3640), .Y (y1607) );
  AO21x1_ASAP7_75t_R   g3868( .A1 (n1838), .A2 (n29), .B (n3867), .Y (y1608) );
  AND2x2_ASAP7_75t_R   g3869( .A (y1393), .B (n455), .Y (y1609) );
  AO33x2_ASAP7_75t_R   g3870( .A1 (n22), .A2 (n672), .A3 (n1838), .B1 (n72), .B2 (n401), .B3 (y2079), .Y (y1610) );
  OR3x1_ASAP7_75t_R    g3871( .A (n529), .B (n962), .C (n12), .Y (n3879) );
  NAND2x1_ASAP7_75t_R  g3872( .A (n12), .B (n1082), .Y (n3880) );
  AND2x2_ASAP7_75t_R   g3873( .A (n3879), .B (n3880), .Y (y1611) );
  AO21x1_ASAP7_75t_R   g3874( .A1 (x0), .A2 (n22), .B (n369), .Y (n3882) );
  AND3x1_ASAP7_75t_R   g3875( .A (n12), .B (n17), .C (x4), .Y (n3883) );
  INVx1_ASAP7_75t_R    g3876( .A (n3883), .Y (n3884) );
  AND2x2_ASAP7_75t_R   g3877( .A (n3882), .B (n3884), .Y (y1612) );
  INVx1_ASAP7_75t_R    g3878( .A (n3218), .Y (y3808) );
  INVx1_ASAP7_75t_R    g3879( .A (n1791), .Y (y2500) );
  AO21x1_ASAP7_75t_R   g3880( .A1 (y3808), .A2 (x0), .B (y2500), .Y (y1613) );
  AND2x2_ASAP7_75t_R   g3881( .A (y432), .B (n556), .Y (y1614) );
  AO21x1_ASAP7_75t_R   g3882( .A1 (n243), .A2 (x0), .B (x2), .Y (n3890) );
  OR3x1_ASAP7_75t_R    g3883( .A (y863), .B (n15), .C (x3), .Y (n3891) );
  INVx1_ASAP7_75t_R    g3884( .A (n3891), .Y (n3892) );
  NOR2x1_ASAP7_75t_R   g3885( .A (n227), .B (n3892), .Y (n3893) );
  OA21x2_ASAP7_75t_R   g3886( .A1 (n3890), .A2 (n261), .B (n3893), .Y (y1615) );
  AO21x1_ASAP7_75t_R   g3887( .A1 (n529), .A2 (n72), .B (n3025), .Y (y1616) );
  AND3x1_ASAP7_75t_R   g3888( .A (n17), .B (n15), .C (x4), .Y (n3896) );
  AO21x1_ASAP7_75t_R   g3889( .A1 (x3), .A2 (x2), .B (n3896), .Y (n3897) );
  OR3x1_ASAP7_75t_R    g3890( .A (n76), .B (y2079), .C (x4), .Y (n3898) );
  INVx1_ASAP7_75t_R    g3891( .A (n3898), .Y (n3899) );
  AO21x1_ASAP7_75t_R   g3892( .A1 (n3897), .A2 (y2079), .B (n3899), .Y (y1617) );
  AO21x1_ASAP7_75t_R   g3893( .A1 (n421), .A2 (n22), .B (x2), .Y (n3901) );
  OR3x1_ASAP7_75t_R    g3894( .A (n756), .B (n17), .C (n22), .Y (n3902) );
  INVx1_ASAP7_75t_R    g3895( .A (n3902), .Y (n3903) );
  AO21x1_ASAP7_75t_R   g3896( .A1 (n3901), .A2 (n382), .B (n3903), .Y (y1618) );
  AO21x1_ASAP7_75t_R   g3897( .A1 (n15), .A2 (x5), .B (x4), .Y (n3905) );
  OR3x1_ASAP7_75t_R    g3898( .A (n164), .B (n163), .C (n3905), .Y (n3906) );
  NAND2x1_ASAP7_75t_R  g3899( .A (x4), .B (n3083), .Y (n3907) );
  AND2x2_ASAP7_75t_R   g3900( .A (n3906), .B (n3907), .Y (y1619) );
  AO21x1_ASAP7_75t_R   g3901( .A1 (n17), .A2 (x5), .B (n15), .Y (n3909) );
  AO32x1_ASAP7_75t_R   g3902( .A1 (x4), .A2 (y2079), .A3 (n72), .B1 (n22), .B2 (n3909), .Y (y1620) );
  NAND2x1_ASAP7_75t_R  g3903( .A (n3480), .B (n1106), .Y (y2305) );
  AND2x2_ASAP7_75t_R   g3904( .A (y2305), .B (n546), .Y (y1621) );
  AO22x1_ASAP7_75t_R   g3905( .A1 (x4), .A2 (y195), .B1 (n22), .B2 (n3696), .Y (y1622) );
  NAND2x1_ASAP7_75t_R  g3906( .A (n15), .B (n3338), .Y (n3914) );
  OA21x2_ASAP7_75t_R   g3907( .A1 (n396), .A2 (n3914), .B (y1287), .Y (y1623) );
  AND3x1_ASAP7_75t_R   g3908( .A (n534), .B (n219), .C (n556), .Y (y1624) );
  AO21x1_ASAP7_75t_R   g3909( .A1 (n3384), .A2 (y2079), .B (n3085), .Y (y1626) );
  AO21x1_ASAP7_75t_R   g3910( .A1 (x2), .A2 (x3), .B (x5), .Y (n3918) );
  NAND2x1_ASAP7_75t_R  g3911( .A (x5), .B (n3024), .Y (n3919) );
  OA21x2_ASAP7_75t_R   g3912( .A1 (n3182), .A2 (n3918), .B (n3919), .Y (y1627) );
  AO21x1_ASAP7_75t_R   g3913( .A1 (n3284), .A2 (x0), .B (n628), .Y (y1628) );
  AO21x1_ASAP7_75t_R   g3914( .A1 (n52), .A2 (n1522), .B (n2839), .Y (n3922) );
  AND2x2_ASAP7_75t_R   g3915( .A (n1515), .B (n3922), .Y (y1629) );
  NAND2x1_ASAP7_75t_R  g3916( .A (x1), .B (n439), .Y (n3924) );
  AND2x2_ASAP7_75t_R   g3917( .A (n3924), .B (n3380), .Y (y1630) );
  OA22x2_ASAP7_75t_R   g3918( .A1 (n22), .A2 (n3005), .B1 (n1163), .B2 (n3004), .Y (y1631) );
  NAND2x1_ASAP7_75t_R  g3919( .A (n856), .B (n290), .Y (n3927) );
  AND3x1_ASAP7_75t_R   g3920( .A (n3927), .B (n3705), .C (n556), .Y (y1632) );
  AND2x2_ASAP7_75t_R   g3921( .A (n290), .B (n360), .Y (n3929) );
  AND2x2_ASAP7_75t_R   g3922( .A (y1693), .B (x2), .Y (n3930) );
  AO21x1_ASAP7_75t_R   g3923( .A1 (n1646), .A2 (n3929), .B (n3930), .Y (y1633) );
  AO21x1_ASAP7_75t_R   g3924( .A1 (n455), .A2 (n43), .B (y767), .Y (y1634) );
  AO21x1_ASAP7_75t_R   g3925( .A1 (n29), .A2 (n1838), .B (n1269), .Y (y1636) );
  AND2x2_ASAP7_75t_R   g3926( .A (n3866), .B (n3025), .Y (n3934) );
  AO21x1_ASAP7_75t_R   g3927( .A1 (n401), .A2 (n1269), .B (n3934), .Y (y1637) );
  NAND2x1_ASAP7_75t_R  g3928( .A (x2), .B (n2256), .Y (n3936) );
  INVx1_ASAP7_75t_R    g3929( .A (n3936), .Y (n3937) );
  OA21x2_ASAP7_75t_R   g3930( .A1 (n3937), .A2 (y863), .B (n1657), .Y (y1638) );
  NAND2x1_ASAP7_75t_R  g3931( .A (n3123), .B (n3469), .Y (n3939) );
  AND2x2_ASAP7_75t_R   g3932( .A (n3939), .B (n17), .Y (n3940) );
  AO21x1_ASAP7_75t_R   g3933( .A1 (n3630), .A2 (x3), .B (n3940), .Y (y1639) );
  OA21x2_ASAP7_75t_R   g3934( .A1 (n1265), .A2 (n1158), .B (y1540), .Y (y1640) );
  AO21x1_ASAP7_75t_R   g3935( .A1 (x5), .A2 (n17), .B (n3567), .Y (n3943) );
  AO21x1_ASAP7_75t_R   g3936( .A1 (y2079), .A2 (x2), .B (n22), .Y (n3944) );
  AND2x2_ASAP7_75t_R   g3937( .A (n3943), .B (n3944), .Y (y1641) );
  NAND2x1_ASAP7_75t_R  g3938( .A (n28), .B (n740), .Y (n3946) );
  AND2x2_ASAP7_75t_R   g3939( .A (n3946), .B (n3705), .Y (y1642) );
  AO21x1_ASAP7_75t_R   g3940( .A1 (n63), .A2 (n64), .B (x3), .Y (n3948) );
  INVx1_ASAP7_75t_R    g3941( .A (n3948), .Y (n3949) );
  AO21x1_ASAP7_75t_R   g3942( .A1 (n125), .A2 (n277), .B (n3949), .Y (y1643) );
  AO21x1_ASAP7_75t_R   g3943( .A1 (n3298), .A2 (x3), .B (n3294), .Y (n3951) );
  XOR2x2_ASAP7_75t_R   g3944( .A (n3951), .B (n22), .Y (y1644) );
  AO221x2_ASAP7_75t_R  g3945( .A1 (n12), .A2 (y2079), .B1 (n700), .B2 (n537), .C (n442), .Y (y1645) );
  AO21x1_ASAP7_75t_R   g3946( .A1 (n29), .A2 (n1838), .B (n3819), .Y (y1646) );
  INVx1_ASAP7_75t_R    g3947( .A (n2169), .Y (n3955) );
  AOI21x1_ASAP7_75t_R  g3948( .A1 (n3955), .A2 (n1841), .B (n1134), .Y (y1647) );
  AND2x2_ASAP7_75t_R   g3949( .A (n2003), .B (n1188), .Y (y1648) );
  AND3x1_ASAP7_75t_R   g3950( .A (y9), .B (n482), .C (n556), .Y (y1649) );
  AND3x1_ASAP7_75t_R   g3951( .A (n1891), .B (n908), .C (n299), .Y (y1650) );
  AND2x2_ASAP7_75t_R   g3952( .A (n137), .B (y2079), .Y (n3960) );
  OA21x2_ASAP7_75t_R   g3953( .A1 (n3960), .A2 (n3025), .B (n3927), .Y (y1651) );
  OA21x2_ASAP7_75t_R   g3954( .A1 (n481), .A2 (n511), .B (n387), .Y (y1652) );
  AND3x1_ASAP7_75t_R   g3955( .A (n137), .B (n72), .C (y2079), .Y (n3963) );
  AO21x1_ASAP7_75t_R   g3956( .A1 (n77), .A2 (n29), .B (n3963), .Y (y1653) );
  NOR2x1_ASAP7_75t_R   g3957( .A (n312), .B (n746), .Y (n3965) );
  INVx1_ASAP7_75t_R    g3958( .A (n3965), .Y (n3966) );
  AND2x2_ASAP7_75t_R   g3959( .A (n3966), .B (n1445), .Y (y1654) );
  AO21x1_ASAP7_75t_R   g3960( .A1 (n1265), .A2 (n3567), .B (n17), .Y (n3968) );
  OA21x2_ASAP7_75t_R   g3961( .A1 (n3960), .A2 (n22), .B (n3968), .Y (y1655) );
  AO21x1_ASAP7_75t_R   g3962( .A1 (n1082), .A2 (x0), .B (n529), .Y (y1656) );
  AO21x1_ASAP7_75t_R   g3963( .A1 (n1564), .A2 (n63), .B (n17), .Y (n3971) );
  AND2x2_ASAP7_75t_R   g3964( .A (n3971), .B (n236), .Y (y1657) );
  AND3x1_ASAP7_75t_R   g3965( .A (y3293), .B (n84), .C (n3832), .Y (y1658) );
  NOR2x1_ASAP7_75t_R   g3966( .A (n25), .B (n23), .Y (n3974) );
  AND2x2_ASAP7_75t_R   g3967( .A (n604), .B (n1082), .Y (y1675) );
  OR3x1_ASAP7_75t_R    g3968( .A (n3974), .B (y2196), .C (y1675), .Y (y1659) );
  NAND2x1_ASAP7_75t_R  g3969( .A (y2466), .B (n84), .Y (n3977) );
  AND3x1_ASAP7_75t_R   g3970( .A (n12), .B (x3), .C (x4), .Y (n3978) );
  INVx1_ASAP7_75t_R    g3971( .A (n3978), .Y (n3979) );
  AND3x1_ASAP7_75t_R   g3972( .A (n3977), .B (y1343), .C (n3979), .Y (y1660) );
  OR3x1_ASAP7_75t_R    g3973( .A (n518), .B (x2), .C (x3), .Y (n3981) );
  OAI21x1_ASAP7_75t_R  g3974( .A1 (x5), .A2 (n3317), .B (n3981), .Y (y1661) );
  AO21x1_ASAP7_75t_R   g3975( .A1 (n17), .A2 (y2079), .B (n756), .Y (n3983) );
  INVx1_ASAP7_75t_R    g3976( .A (n3983), .Y (n3984) );
  OA21x2_ASAP7_75t_R   g3977( .A1 (n3984), .A2 (n163), .B (n2998), .Y (y1662) );
  AND3x1_ASAP7_75t_R   g3978( .A (n218), .B (y2079), .C (n22), .Y (y1802) );
  INVx1_ASAP7_75t_R    g3979( .A (y1802), .Y (n3987) );
  NAND2x1_ASAP7_75t_R  g3980( .A (x5), .B (n3134), .Y (y3831) );
  AND3x1_ASAP7_75t_R   g3981( .A (n137), .B (n72), .C (x4), .Y (n3989) );
  INVx1_ASAP7_75t_R    g3982( .A (n3989), .Y (n3990) );
  AND3x1_ASAP7_75t_R   g3983( .A (n3987), .B (y3831), .C (n3990), .Y (y1663) );
  AND3x1_ASAP7_75t_R   g3984( .A (n137), .B (n72), .C (n22), .Y (n3992) );
  NAND2x1_ASAP7_75t_R  g3985( .A (y2079), .B (n3992), .Y (n3993) );
  AND2x2_ASAP7_75t_R   g3986( .A (n3993), .B (n556), .Y (y1664) );
  AO21x1_ASAP7_75t_R   g3987( .A1 (n3124), .A2 (n1838), .B (n3611), .Y (y1665) );
  AO21x1_ASAP7_75t_R   g3988( .A1 (n489), .A2 (n490), .B (n503), .Y (y1666) );
  AND2x2_ASAP7_75t_R   g3989( .A (n2478), .B (n219), .Y (n3997) );
  OA21x2_ASAP7_75t_R   g3990( .A1 (n3997), .A2 (x4), .B (n718), .Y (y1667) );
  AO21x1_ASAP7_75t_R   g3991( .A1 (n143), .A2 (x2), .B (x3), .Y (n3999) );
  INVx1_ASAP7_75t_R    g3992( .A (n3999), .Y (n4000) );
  AO21x1_ASAP7_75t_R   g3993( .A1 (n2757), .A2 (n1564), .B (n4000), .Y (y1668) );
  AND2x2_ASAP7_75t_R   g3994( .A (y1777), .B (n632), .Y (y1669) );
  AND2x2_ASAP7_75t_R   g3995( .A (n2720), .B (n2721), .Y (y1670) );
  AND2x2_ASAP7_75t_R   g3996( .A (y1693), .B (n661), .Y (y1671) );
  NAND2x1_ASAP7_75t_R  g3997( .A (n15), .B (n258), .Y (n4005) );
  AO21x1_ASAP7_75t_R   g3998( .A1 (n90), .A2 (n219), .B (n45), .Y (n4006) );
  OA21x2_ASAP7_75t_R   g3999( .A1 (n221), .A2 (n4005), .B (n4006), .Y (y1672) );
  AO21x1_ASAP7_75t_R   g4000( .A1 (n3794), .A2 (n3316), .B (n3132), .Y (y1673) );
  INVx1_ASAP7_75t_R    g4001( .A (n3828), .Y (n4009) );
  AND3x1_ASAP7_75t_R   g4002( .A (n97), .B (n740), .C (x3), .Y (n4010) );
  INVx1_ASAP7_75t_R    g4003( .A (n4010), .Y (n4011) );
  OA21x2_ASAP7_75t_R   g4004( .A1 (n4009), .A2 (n3626), .B (n4011), .Y (y1674) );
  AO21x1_ASAP7_75t_R   g4005( .A1 (n3819), .A2 (x3), .B (n3316), .Y (y1676) );
  AO21x1_ASAP7_75t_R   g4006( .A1 (n12), .A2 (x5), .B (x3), .Y (n4014) );
  NOR2x1_ASAP7_75t_R   g4007( .A (x4), .B (n4014), .Y (n4015) );
  INVx1_ASAP7_75t_R    g4008( .A (n4015), .Y (n4016) );
  AND2x2_ASAP7_75t_R   g4009( .A (y1903), .B (n4016), .Y (y1677) );
  NAND2x1_ASAP7_75t_R  g4010( .A (x2), .B (n3443), .Y (n4018) );
  INVx1_ASAP7_75t_R    g4011( .A (n4018), .Y (n4019) );
  AO21x1_ASAP7_75t_R   g4012( .A1 (n1838), .A2 (n3124), .B (n4019), .Y (y1678) );
  AO21x1_ASAP7_75t_R   g4013( .A1 (x1), .A2 (n22), .B (n538), .Y (y1679) );
  AO21x1_ASAP7_75t_R   g4014( .A1 (n17), .A2 (x5), .B (x2), .Y (n4022) );
  AND2x2_ASAP7_75t_R   g4015( .A (n3302), .B (n4022), .Y (y1680) );
  OR3x1_ASAP7_75t_R    g4016( .A (n81), .B (x5), .C (x4), .Y (n4024) );
  AND2x2_ASAP7_75t_R   g4017( .A (y2016), .B (n4024), .Y (y1681) );
  AO21x1_ASAP7_75t_R   g4018( .A1 (n16), .A2 (n2276), .B (n1208), .Y (n4026) );
  INVx1_ASAP7_75t_R    g4019( .A (n4026), .Y (y1682) );
  INVx1_ASAP7_75t_R    g4020( .A (n3480), .Y (n4028) );
  AO21x1_ASAP7_75t_R   g4021( .A1 (n4028), .A2 (n312), .B (n1907), .Y (y1683) );
  AND3x1_ASAP7_75t_R   g4022( .A (n2999), .B (y2079), .C (n17), .Y (n4030) );
  INVx1_ASAP7_75t_R    g4023( .A (n4030), .Y (n4031) );
  AND3x1_ASAP7_75t_R   g4024( .A (n4031), .B (n3835), .C (y3293), .Y (y1684) );
  AO21x1_ASAP7_75t_R   g4025( .A1 (n15), .A2 (n22), .B (x5), .Y (n4033) );
  AND2x2_ASAP7_75t_R   g4026( .A (n28), .B (n4033), .Y (n4034) );
  INVx1_ASAP7_75t_R    g4027( .A (n4034), .Y (n4035) );
  AND2x2_ASAP7_75t_R   g4028( .A (n4035), .B (n3835), .Y (y1685) );
  NAND2x1_ASAP7_75t_R  g4029( .A (x3), .B (n3823), .Y (n4037) );
  AND3x1_ASAP7_75t_R   g4030( .A (y2079), .B (n22), .C (x2), .Y (n4038) );
  INVx1_ASAP7_75t_R    g4031( .A (n4038), .Y (n4039) );
  AO32x1_ASAP7_75t_R   g4032( .A1 (y3293), .A2 (n4037), .A3 (n4039), .B1 (n1269), .B2 (n1158), .Y (y1686) );
  NAND2x1_ASAP7_75t_R  g4033( .A (n180), .B (n56), .Y (y1687) );
  NOR2x1_ASAP7_75t_R   g4034( .A (x4), .B (n3285), .Y (n4042) );
  OR3x1_ASAP7_75t_R    g4035( .A (n4042), .B (n3294), .C (n529), .Y (y1688) );
  AND2x2_ASAP7_75t_R   g4036( .A (n1275), .B (n1188), .Y (y1689) );
  AO21x1_ASAP7_75t_R   g4037( .A1 (x5), .A2 (n1150), .B (n529), .Y (y1690) );
  AO21x1_ASAP7_75t_R   g4038( .A1 (y1378), .A2 (n17), .B (n959), .Y (y1691) );
  INVx1_ASAP7_75t_R    g4039( .A (n430), .Y (n4047) );
  INVx1_ASAP7_75t_R    g4040( .A (n607), .Y (n4048) );
  OA33x2_ASAP7_75t_R   g4041( .A1 (n16), .A2 (n4047), .A3 (n3149), .B1 (x1), .B2 (n29), .B3 (n4048), .Y (y1692) );
  NAND2x1_ASAP7_75t_R  g4042( .A (n17), .B (n3780), .Y (n4050) );
  OAI21x1_ASAP7_75t_R  g4043( .A1 (n17), .A2 (n4034), .B (n4050), .Y (y1694) );
  AO21x1_ASAP7_75t_R   g4044( .A1 (x5), .A2 (x4), .B (n211), .Y (n4052) );
  NOR2x1_ASAP7_75t_R   g4045( .A (n4052), .B (n4030), .Y (y1695) );
  AND2x2_ASAP7_75t_R   g4046( .A (y802), .B (n228), .Y (y1696) );
  AND3x1_ASAP7_75t_R   g4047( .A (n15), .B (n22), .C (x5), .Y (n4055) );
  INVx1_ASAP7_75t_R    g4048( .A (n4055), .Y (n4056) );
  AO21x1_ASAP7_75t_R   g4049( .A1 (y2079), .A2 (x2), .B (n4055), .Y (n4057) );
  AO32x1_ASAP7_75t_R   g4050( .A1 (n17), .A2 (n4056), .A3 (n3028), .B1 (x3), .B2 (n4057), .Y (y1697) );
  AO21x1_ASAP7_75t_R   g4051( .A1 (n3013), .A2 (n3011), .B (n17), .Y (n4059) );
  OA21x2_ASAP7_75t_R   g4052( .A1 (n3012), .A2 (n391), .B (n4059), .Y (y1698) );
  INVx1_ASAP7_75t_R    g4053( .A (n367), .Y (n4061) );
  AND3x1_ASAP7_75t_R   g4054( .A (n378), .B (y2079), .C (x2), .Y (n4062) );
  NOR2x1_ASAP7_75t_R   g4055( .A (n4061), .B (n4062), .Y (y1699) );
  AND2x2_ASAP7_75t_R   g4056( .A (n3977), .B (y1343), .Y (y1700) );
  AO21x1_ASAP7_75t_R   g4057( .A1 (n1851), .A2 (y2079), .B (n3338), .Y (n4065) );
  AND2x2_ASAP7_75t_R   g4058( .A (n4065), .B (n1620), .Y (y1701) );
  AO21x1_ASAP7_75t_R   g4059( .A1 (y2079), .A2 (x0), .B (n337), .Y (y1702) );
  AND2x2_ASAP7_75t_R   g4060( .A (n185), .B (y2079), .Y (n4068) );
  OR3x1_ASAP7_75t_R    g4061( .A (n1541), .B (n262), .C (n4068), .Y (y1703) );
  OR3x1_ASAP7_75t_R    g4062( .A (x3), .B (x2), .C (x4), .Y (n4070) );
  AND2x2_ASAP7_75t_R   g4063( .A (y1359), .B (n4070), .Y (y1704) );
  AO21x1_ASAP7_75t_R   g4064( .A1 (n3156), .A2 (y2079), .B (y2259), .Y (y1705) );
  AO32x1_ASAP7_75t_R   g4065( .A1 (n360), .A2 (n290), .A3 (n3662), .B1 (n378), .B2 (n3661), .Y (y1706) );
  AND2x2_ASAP7_75t_R   g4066( .A (y232), .B (n1510), .Y (y1707) );
  INVx1_ASAP7_75t_R    g4067( .A (n3284), .Y (n4075) );
  AO21x1_ASAP7_75t_R   g4068( .A1 (n319), .A2 (x4), .B (n3285), .Y (n4076) );
  INVx1_ASAP7_75t_R    g4069( .A (n4076), .Y (n4077) );
  AO21x1_ASAP7_75t_R   g4070( .A1 (n3285), .A2 (n4075), .B (n4077), .Y (n4078) );
  AO21x1_ASAP7_75t_R   g4071( .A1 (n15), .A2 (y2079), .B (n4078), .Y (y1708) );
  INVx1_ASAP7_75t_R    g4072( .A (n926), .Y (y1709) );
  INVx1_ASAP7_75t_R    g4073( .A (n3766), .Y (n4081) );
  AO21x1_ASAP7_75t_R   g4074( .A1 (n1050), .A2 (n1743), .B (n4081), .Y (n4082) );
  OR3x1_ASAP7_75t_R    g4075( .A (y2466), .B (n12), .C (x1), .Y (n4083) );
  AND2x2_ASAP7_75t_R   g4076( .A (n4082), .B (n4083), .Y (y1710) );
  AND2x2_ASAP7_75t_R   g4077( .A (n1923), .B (n1188), .Y (n4085) );
  NOR2x1_ASAP7_75t_R   g4078( .A (x5), .B (n4085), .Y (n4086) );
  AO21x1_ASAP7_75t_R   g4079( .A1 (x5), .A2 (n914), .B (n4086), .Y (y1711) );
  AND3x1_ASAP7_75t_R   g4080( .A (x3), .B (x2), .C (x5), .Y (n4088) );
  INVx1_ASAP7_75t_R    g4081( .A (n4088), .Y (n4089) );
  AO21x1_ASAP7_75t_R   g4082( .A1 (n4089), .A2 (n1572), .B (n22), .Y (n4090) );
  AND2x2_ASAP7_75t_R   g4083( .A (n4090), .B (n3134), .Y (y1712) );
  AND2x2_ASAP7_75t_R   g4084( .A (n3987), .B (y3831), .Y (y1713) );
  AO21x1_ASAP7_75t_R   g4085( .A1 (y1356), .A2 (x2), .B (n2126), .Y (y1715) );
  AND3x1_ASAP7_75t_R   g4086( .A (n360), .B (n3469), .C (x5), .Y (n4094) );
  NOR2x1_ASAP7_75t_R   g4087( .A (n164), .B (n4094), .Y (y1716) );
  AO21x1_ASAP7_75t_R   g4088( .A1 (y9), .A2 (n211), .B (n143), .Y (n4096) );
  AO21x1_ASAP7_75t_R   g4089( .A1 (n2556), .A2 (n16), .B (n4096), .Y (y1717) );
  AO21x1_ASAP7_75t_R   g4090( .A1 (n1693), .A2 (n258), .B (n2419), .Y (y1718) );
  AO21x1_ASAP7_75t_R   g4091( .A1 (n22), .A2 (y2079), .B (n17), .Y (n4099) );
  INVx1_ASAP7_75t_R    g4092( .A (n4099), .Y (n4100) );
  NOR2x1_ASAP7_75t_R   g4093( .A (x4), .B (x2), .Y (n4101) );
  INVx1_ASAP7_75t_R    g4094( .A (n3804), .Y (n4102) );
  AO21x1_ASAP7_75t_R   g4095( .A1 (n369), .A2 (n4101), .B (n4102), .Y (n4103) );
  AOI22x1_ASAP7_75t_R  g4096( .A1 (x2), .A2 (n4100), .B1 (n4103), .B2 (x5), .Y (y1719) );
  OR3x1_ASAP7_75t_R    g4097( .A (n3203), .B (n484), .C (n527), .Y (n4105) );
  AND2x2_ASAP7_75t_R   g4098( .A (n4105), .B (y250), .Y (y1720) );
  AO21x1_ASAP7_75t_R   g4099( .A1 (n15), .A2 (n17), .B (x4), .Y (n4107) );
  NAND2x1_ASAP7_75t_R  g4100( .A (x5), .B (n4107), .Y (n4108) );
  AO21x1_ASAP7_75t_R   g4101( .A1 (x5), .A2 (n15), .B (n360), .Y (n4109) );
  AND2x2_ASAP7_75t_R   g4102( .A (n4108), .B (n4109), .Y (y1721) );
  OR3x1_ASAP7_75t_R    g4103( .A (n3203), .B (x5), .C (x3), .Y (n4111) );
  OA21x2_ASAP7_75t_R   g4104( .A1 (n671), .A2 (y1702), .B (n4111), .Y (y1722) );
  OR3x1_ASAP7_75t_R    g4105( .A (n2099), .B (n271), .C (n262), .Y (y1723) );
  AND2x2_ASAP7_75t_R   g4106( .A (n218), .B (n29), .Y (n4114) );
  OR3x1_ASAP7_75t_R    g4107( .A (n4114), .B (n3132), .C (n3896), .Y (y1724) );
  INVx1_ASAP7_75t_R    g4108( .A (n4014), .Y (n4116) );
  AO21x1_ASAP7_75t_R   g4109( .A1 (n12), .A2 (n17), .B (x4), .Y (n4117) );
  AO21x1_ASAP7_75t_R   g4110( .A1 (y3852), .A2 (x3), .B (n4117), .Y (n4118) );
  OA21x2_ASAP7_75t_R   g4111( .A1 (n4116), .A2 (n718), .B (n4118), .Y (y1725) );
  OAI21x1_ASAP7_75t_R  g4112( .A1 (n2715), .A2 (n1051), .B (n1111), .Y (y1726) );
  AO21x1_ASAP7_75t_R   g4113( .A1 (n12), .A2 (n961), .B (n1132), .Y (y1727) );
  AND2x2_ASAP7_75t_R   g4114( .A (n556), .B (n1047), .Y (n4122) );
  AO21x1_ASAP7_75t_R   g4115( .A1 (n4122), .A2 (n534), .B (n2001), .Y (y1728) );
  INVx1_ASAP7_75t_R    g4116( .A (n4107), .Y (n4124) );
  AO21x1_ASAP7_75t_R   g4117( .A1 (n4124), .A2 (n3828), .B (n529), .Y (y1729) );
  AO21x1_ASAP7_75t_R   g4118( .A1 (n218), .A2 (n29), .B (n529), .Y (y1730) );
  AO21x1_ASAP7_75t_R   g4119( .A1 (n466), .A2 (n58), .B (n1775), .Y (y1731) );
  OA21x2_ASAP7_75t_R   g4120( .A1 (n2551), .A2 (n145), .B (n2552), .Y (y1732) );
  INVx1_ASAP7_75t_R    g4121( .A (n3310), .Y (n4129) );
  AO21x1_ASAP7_75t_R   g4122( .A1 (n4129), .A2 (n348), .B (y2079), .Y (n4130) );
  OAI21x1_ASAP7_75t_R  g4123( .A1 (n3310), .A2 (n285), .B (n4130), .Y (n4131) );
  AO21x1_ASAP7_75t_R   g4124( .A1 (x2), .A2 (n382), .B (n4131), .Y (y1733) );
  AO21x1_ASAP7_75t_R   g4125( .A1 (n740), .A2 (n43), .B (y773), .Y (y1734) );
  AO21x1_ASAP7_75t_R   g4126( .A1 (n474), .A2 (n1059), .B (n529), .Y (y1735) );
  NAND2x1_ASAP7_75t_R  g4127( .A (n292), .B (n290), .Y (y3132) );
  INVx1_ASAP7_75t_R    g4128( .A (y3132), .Y (n4136) );
  AND2x2_ASAP7_75t_R   g4129( .A (y3132), .B (x2), .Y (n4137) );
  AO21x1_ASAP7_75t_R   g4130( .A1 (n15), .A2 (n4136), .B (n4137), .Y (y1736) );
  INVx1_ASAP7_75t_R    g4131( .A (n459), .Y (n4139) );
  AO21x1_ASAP7_75t_R   g4132( .A1 (n1370), .A2 (y1894), .B (n4139), .Y (y1737) );
  AND3x1_ASAP7_75t_R   g4133( .A (y9), .B (n1453), .C (y2079), .Y (y1738) );
  OR3x1_ASAP7_75t_R    g4134( .A (y2466), .B (x2), .C (x3), .Y (n4142) );
  AND2x2_ASAP7_75t_R   g4135( .A (n4142), .B (y1359), .Y (y1739) );
  AND2x2_ASAP7_75t_R   g4136( .A (n2276), .B (n883), .Y (y1740) );
  AO21x1_ASAP7_75t_R   g4137( .A1 (n174), .A2 (n1312), .B (n262), .Y (y1741) );
  AO21x1_ASAP7_75t_R   g4138( .A1 (y2079), .A2 (x3), .B (n638), .Y (y1742) );
  AND2x2_ASAP7_75t_R   g4139( .A (y1359), .B (n1572), .Y (y1743) );
  AO21x1_ASAP7_75t_R   g4140( .A1 (y2079), .A2 (n174), .B (n272), .Y (y1744) );
  NAND2x1_ASAP7_75t_R  g4141( .A (n22), .B (n3828), .Y (n4149) );
  INVx1_ASAP7_75t_R    g4142( .A (n4149), .Y (n4150) );
  OR3x1_ASAP7_75t_R    g4143( .A (y2466), .B (x3), .C (x2), .Y (n4151) );
  OA21x2_ASAP7_75t_R   g4144( .A1 (n4150), .A2 (n3774), .B (n4151), .Y (y1745) );
  AO21x1_ASAP7_75t_R   g4145( .A1 (y2079), .A2 (n348), .B (n3189), .Y (y2900) );
  AND2x2_ASAP7_75t_R   g4146( .A (y2900), .B (n382), .Y (y1746) );
  AO21x1_ASAP7_75t_R   g4147( .A1 (n12), .A2 (n28), .B (n300), .Y (n4155) );
  AO221x2_ASAP7_75t_R  g4148( .A1 (x1), .A2 (n23), .B1 (n16), .B2 (n4155), .C (n529), .Y (y1747) );
  AND2x2_ASAP7_75t_R   g4149( .A (y3198), .B (n3797), .Y (y1748) );
  AND3x1_ASAP7_75t_R   g4150( .A (n2298), .B (n1490), .C (y2079), .Y (y1749) );
  AO21x1_ASAP7_75t_R   g4151( .A1 (y1356), .A2 (x2), .B (n2178), .Y (y1750) );
  AND3x1_ASAP7_75t_R   g4152( .A (y3377), .B (n724), .C (x0), .Y (y1752) );
  AO32x1_ASAP7_75t_R   g4153( .A1 (n299), .A2 (x3), .A3 (y2079), .B1 (n604), .B2 (n3116), .Y (y1753) );
  AO21x1_ASAP7_75t_R   g4154( .A1 (n671), .A2 (n22), .B (x0), .Y (n4162) );
  AND2x2_ASAP7_75t_R   g4155( .A (n600), .B (n4162), .Y (y1754) );
  AO32x1_ASAP7_75t_R   g4156( .A1 (n22), .A2 (n3089), .A3 (n3579), .B1 (x0), .B2 (n3443), .Y (y1755) );
  OR3x1_ASAP7_75t_R    g4157( .A (n418), .B (n16), .C (n12), .Y (n4165) );
  INVx1_ASAP7_75t_R    g4158( .A (n4165), .Y (n4166) );
  AO21x1_ASAP7_75t_R   g4159( .A1 (n1223), .A2 (n3148), .B (n4166), .Y (n4167) );
  AND2x2_ASAP7_75t_R   g4160( .A (n4167), .B (y3293), .Y (y1756) );
  AND2x2_ASAP7_75t_R   g4161( .A (y3293), .B (y1894), .Y (y1757) );
  AND3x1_ASAP7_75t_R   g4162( .A (n556), .B (n77), .C (n4070), .Y (y1758) );
  OR3x1_ASAP7_75t_R    g4163( .A (n756), .B (x4), .C (x3), .Y (n4171) );
  AND3x1_ASAP7_75t_R   g4164( .A (n4011), .B (n4171), .C (n556), .Y (y1759) );
  AO21x1_ASAP7_75t_R   g4165( .A1 (n455), .A2 (n765), .B (n437), .Y (n4173) );
  AND3x1_ASAP7_75t_R   g4166( .A (n4173), .B (n2940), .C (n299), .Y (y1760) );
  NOR2x1_ASAP7_75t_R   g4167( .A (x3), .B (n429), .Y (n4175) );
  NOR2x1_ASAP7_75t_R   g4168( .A (n3598), .B (n4175), .Y (y1761) );
  AO21x1_ASAP7_75t_R   g4169( .A1 (y2079), .A2 (n125), .B (n3386), .Y (y2034) );
  AND2x2_ASAP7_75t_R   g4170( .A (y2034), .B (n84), .Y (y1763) );
  OA211x2_ASAP7_75t_R  g4171( .A1 (x0), .A2 (n1190), .B (n919), .C (n455), .Y (y1764) );
  AND3x1_ASAP7_75t_R   g4172( .A (n17), .B (y2079), .C (x2), .Y (n4180) );
  NOR2x1_ASAP7_75t_R   g4173( .A (n4180), .B (n407), .Y (y1765) );
  OA22x2_ASAP7_75t_R   g4174( .A1 (n16), .A2 (n2493), .B1 (x1), .B2 (n2137), .Y (y1766) );
  AO21x1_ASAP7_75t_R   g4175( .A1 (n3443), .A2 (x0), .B (n337), .Y (y1767) );
  AO32x1_ASAP7_75t_R   g4176( .A1 (n22), .A2 (n583), .A3 (n2180), .B1 (n971), .B2 (n908), .Y (y1768) );
  AND3x1_ASAP7_75t_R   g4177( .A (n369), .B (n290), .C (x0), .Y (y1793) );
  AO21x1_ASAP7_75t_R   g4178( .A1 (n12), .A2 (n641), .B (y1793), .Y (y1769) );
  AO32x1_ASAP7_75t_R   g4179( .A1 (y3293), .A2 (n1222), .A3 (n3148), .B1 (y2079), .B2 (n3450), .Y (y1770) );
  AO21x1_ASAP7_75t_R   g4180( .A1 (y2079), .A2 (x2), .B (n347), .Y (n4188) );
  INVx1_ASAP7_75t_R    g4181( .A (n4188), .Y (n4189) );
  AND3x1_ASAP7_75t_R   g4182( .A (n360), .B (n97), .C (n290), .Y (n4190) );
  NOR2x1_ASAP7_75t_R   g4183( .A (n4189), .B (n4190), .Y (y1771) );
  INVx1_ASAP7_75t_R    g4184( .A (y2813), .Y (n4192) );
  OA331x2_ASAP7_75t_R  g4185( .A1 (x2), .A2 (n3487), .A3 (n4192), .B1 (n15), .B2 (y2079), .B3 (y863), .C1 (n228), .Y (y1772) );
  AND3x1_ASAP7_75t_R   g4186( .A (n1265), .B (n137), .C (n406), .Y (y1773) );
  AO21x1_ASAP7_75t_R   g4187( .A1 (y2079), .A2 (n360), .B (n3009), .Y (n4195) );
  AO21x1_ASAP7_75t_R   g4188( .A1 (n537), .A2 (n17), .B (n4195), .Y (y1774) );
  AND2x2_ASAP7_75t_R   g4189( .A (n84), .B (n125), .Y (n4197) );
  OA21x2_ASAP7_75t_R   g4190( .A1 (n4197), .A2 (x5), .B (y3198), .Y (y1776) );
  NAND2x1_ASAP7_75t_R  g4191( .A (n740), .B (n1467), .Y (y1778) );
  AO21x1_ASAP7_75t_R   g4192( .A1 (x3), .A2 (x2), .B (y2079), .Y (n4200) );
  AO21x1_ASAP7_75t_R   g4193( .A1 (n22), .A2 (n4200), .B (n3132), .Y (n4201) );
  NOR2x1_ASAP7_75t_R   g4194( .A (n3567), .B (n316), .Y (n4202) );
  INVx1_ASAP7_75t_R    g4195( .A (n4202), .Y (n4203) );
  OA21x2_ASAP7_75t_R   g4196( .A1 (n81), .A2 (n4201), .B (n4203), .Y (y1779) );
  AO21x1_ASAP7_75t_R   g4197( .A1 (n22), .A2 (x5), .B (n145), .Y (n4205) );
  OA21x2_ASAP7_75t_R   g4198( .A1 (n4205), .A2 (n315), .B (n3327), .Y (y1780) );
  AND3x1_ASAP7_75t_R   g4199( .A (n1114), .B (n453), .C (y3852), .Y (y1781) );
  AND3x1_ASAP7_75t_R   g4200( .A (n451), .B (n3979), .C (y1281), .Y (y1782) );
  INVx1_ASAP7_75t_R    g4201( .A (n192), .Y (n4209) );
  AO21x1_ASAP7_75t_R   g4202( .A1 (n4209), .A2 (y263), .B (n214), .Y (y1783) );
  AO21x1_ASAP7_75t_R   g4203( .A1 (n63), .A2 (n851), .B (x3), .Y (n4211) );
  AO21x1_ASAP7_75t_R   g4204( .A1 (n90), .A2 (n15), .B (n2731), .Y (n4212) );
  AND2x2_ASAP7_75t_R   g4205( .A (n4211), .B (n4212), .Y (n4213) );
  AOI21x1_ASAP7_75t_R  g4206( .A1 (n12), .A2 (n129), .B (n4213), .Y (y1784) );
  AND3x1_ASAP7_75t_R   g4207( .A (n455), .B (n463), .C (x0), .Y (y1785) );
  AO21x1_ASAP7_75t_R   g4208( .A1 (n15), .A2 (x5), .B (x3), .Y (n4216) );
  NOR2x1_ASAP7_75t_R   g4209( .A (x4), .B (n4216), .Y (n4217) );
  NOR2x1_ASAP7_75t_R   g4210( .A (n3118), .B (n4217), .Y (y1786) );
  AND2x2_ASAP7_75t_R   g4211( .A (n455), .B (n219), .Y (n4219) );
  AO21x1_ASAP7_75t_R   g4212( .A1 (n4219), .A2 (n1191), .B (n532), .Y (y1787) );
  AND3x1_ASAP7_75t_R   g4213( .A (n2323), .B (n2509), .C (n219), .Y (y1788) );
  OA22x2_ASAP7_75t_R   g4214( .A1 (n1319), .A2 (n3105), .B1 (y1456), .B2 (n644), .Y (y1789) );
  AO21x1_ASAP7_75t_R   g4215( .A1 (y2079), .A2 (n3989), .B (n3135), .Y (y1790) );
  AO21x1_ASAP7_75t_R   g4216( .A1 (n1305), .A2 (x2), .B (n1380), .Y (y1791) );
  INVx1_ASAP7_75t_R    g4217( .A (n3040), .Y (n4225) );
  AND3x1_ASAP7_75t_R   g4218( .A (n369), .B (n360), .C (n290), .Y (y2740) );
  AO21x1_ASAP7_75t_R   g4219( .A1 (x5), .A2 (n4225), .B (y2740), .Y (y1792) );
  OR3x1_ASAP7_75t_R    g4220( .A (n418), .B (n17), .C (x0), .Y (n4228) );
  AND2x2_ASAP7_75t_R   g4221( .A (n615), .B (n4228), .Y (y1794) );
  AND3x1_ASAP7_75t_R   g4222( .A (n672), .B (n1838), .C (n22), .Y (n4230) );
  AO21x1_ASAP7_75t_R   g4223( .A1 (y2079), .A2 (x2), .B (n4230), .Y (y1795) );
  OR3x1_ASAP7_75t_R    g4224( .A (x2), .B (x4), .C (x3), .Y (n4232) );
  AO21x1_ASAP7_75t_R   g4225( .A1 (n22), .A2 (n17), .B (n15), .Y (n4233) );
  NAND2x1_ASAP7_75t_R  g4226( .A (n4232), .B (n4233), .Y (n4234) );
  OR3x1_ASAP7_75t_R    g4227( .A (n347), .B (y2079), .C (n15), .Y (n4235) );
  OA21x2_ASAP7_75t_R   g4228( .A1 (n4234), .A2 (n288), .B (n4235), .Y (y1796) );
  AO21x1_ASAP7_75t_R   g4229( .A1 (n28), .A2 (n45), .B (n3298), .Y (y1797) );
  AO21x1_ASAP7_75t_R   g4230( .A1 (x3), .A2 (x4), .B (n756), .Y (n4238) );
  AO21x1_ASAP7_75t_R   g4231( .A1 (n671), .A2 (n22), .B (n4238), .Y (n4239) );
  AND3x1_ASAP7_75t_R   g4232( .A (n756), .B (x4), .C (x3), .Y (n4240) );
  INVx1_ASAP7_75t_R    g4233( .A (n4240), .Y (n4241) );
  AND2x2_ASAP7_75t_R   g4234( .A (n4239), .B (n4241), .Y (y1798) );
  AND2x2_ASAP7_75t_R   g4235( .A (n2971), .B (x4), .Y (n4243) );
  AO21x1_ASAP7_75t_R   g4236( .A1 (n1572), .A2 (n29), .B (n4243), .Y (y1799) );
  AO221x2_ASAP7_75t_R  g4237( .A1 (n537), .A2 (n700), .B1 (n22), .B2 (n997), .C (n363), .Y (y1800) );
  AO21x1_ASAP7_75t_R   g4238( .A1 (y2079), .A2 (x0), .B (n347), .Y (n4246) );
  AND3x1_ASAP7_75t_R   g4239( .A (n3109), .B (n4246), .C (y3176), .Y (y1801) );
  AND2x2_ASAP7_75t_R   g4240( .A (n380), .B (y3176), .Y (y1803) );
  AO21x1_ASAP7_75t_R   g4241( .A1 (x3), .A2 (x5), .B (x4), .Y (n4249) );
  INVx1_ASAP7_75t_R    g4242( .A (n4249), .Y (n4250) );
  AO21x1_ASAP7_75t_R   g4243( .A1 (n84), .A2 (y2079), .B (n4250), .Y (y2238) );
  AND2x2_ASAP7_75t_R   g4244( .A (n1161), .B (y2238), .Y (y1804) );
  AO21x1_ASAP7_75t_R   g4245( .A1 (n1295), .A2 (n1296), .B (n15), .Y (n4253) );
  AO21x1_ASAP7_75t_R   g4246( .A1 (x1), .A2 (n17), .B (n746), .Y (n4254) );
  AND3x1_ASAP7_75t_R   g4247( .A (n4253), .B (n4254), .C (n1480), .Y (y1805) );
  OA21x2_ASAP7_75t_R   g4248( .A1 (n1646), .A2 (n3471), .B (n556), .Y (y1806) );
  AO21x1_ASAP7_75t_R   g4249( .A1 (n1232), .A2 (n2407), .B (y2093), .Y (y1807) );
  AO21x1_ASAP7_75t_R   g4250( .A1 (n401), .A2 (n1269), .B (n3525), .Y (y1808) );
  NAND2x1_ASAP7_75t_R  g4251( .A (n12), .B (n1839), .Y (n4259) );
  AND2x2_ASAP7_75t_R   g4252( .A (n4259), .B (n1838), .Y (n4260) );
  AO21x1_ASAP7_75t_R   g4253( .A1 (n137), .A2 (n72), .B (n16), .Y (n4261) );
  NOR2x1_ASAP7_75t_R   g4254( .A (n12), .B (n4261), .Y (n4262) );
  INVx1_ASAP7_75t_R    g4255( .A (n4262), .Y (n4263) );
  OA21x2_ASAP7_75t_R   g4256( .A1 (y2220), .A2 (n4260), .B (n4263), .Y (y1809) );
  AO21x1_ASAP7_75t_R   g4257( .A1 (x1), .A2 (y2079), .B (n572), .Y (n4265) );
  AND3x1_ASAP7_75t_R   g4258( .A (n4265), .B (n546), .C (y3852), .Y (y1810) );
  AND2x2_ASAP7_75t_R   g4259( .A (n290), .B (n3327), .Y (y1811) );
  AND2x2_ASAP7_75t_R   g4260( .A (y2723), .B (x0), .Y (y1812) );
  INVx1_ASAP7_75t_R    g4261( .A (n718), .Y (n4269) );
  NAND2x1_ASAP7_75t_R  g4262( .A (x3), .B (n4269), .Y (n4270) );
  OA21x2_ASAP7_75t_R   g4263( .A1 (n3172), .A2 (n2843), .B (n4270), .Y (y1813) );
  AND2x2_ASAP7_75t_R   g4264( .A (y2852), .B (n451), .Y (y1814) );
  INVx1_ASAP7_75t_R    g4265( .A (n3285), .Y (n4273) );
  AND3x1_ASAP7_75t_R   g4266( .A (n4273), .B (n290), .C (n28), .Y (n4274) );
  INVx1_ASAP7_75t_R    g4267( .A (n4274), .Y (n4275) );
  AO21x1_ASAP7_75t_R   g4268( .A1 (n28), .A2 (n290), .B (x2), .Y (n4276) );
  AND2x2_ASAP7_75t_R   g4269( .A (n4275), .B (n4276), .Y (y1815) );
  OA22x2_ASAP7_75t_R   g4270( .A1 (n537), .A2 (n463), .B1 (n3450), .B2 (n1980), .Y (y1816) );
  INVx1_ASAP7_75t_R    g4271( .A (n2980), .Y (n4279) );
  NAND2x1_ASAP7_75t_R  g4272( .A (y3377), .B (n4279), .Y (n4280) );
  AND2x2_ASAP7_75t_R   g4273( .A (n4280), .B (n3030), .Y (y1817) );
  NOR2x1_ASAP7_75t_R   g4274( .A (n22), .B (n58), .Y (n4282) );
  OAI22x1_ASAP7_75t_R  g4275( .A1 (n1927), .A2 (n17), .B1 (n4282), .B2 (n3267), .Y (y1818) );
  AO21x1_ASAP7_75t_R   g4276( .A1 (n2315), .A2 (n64), .B (n1339), .Y (y1819) );
  NOR2x1_ASAP7_75t_R   g4277( .A (n756), .B (n4250), .Y (n4285) );
  AND3x1_ASAP7_75t_R   g4278( .A (n756), .B (n22), .C (n17), .Y (n4286) );
  OA21x2_ASAP7_75t_R   g4279( .A1 (n4285), .A2 (n4286), .B (n3469), .Y (y1820) );
  AND3x1_ASAP7_75t_R   g4280( .A (x0), .B (x3), .C (x4), .Y (n4288) );
  INVx1_ASAP7_75t_R    g4281( .A (n4288), .Y (n4289) );
  AND2x2_ASAP7_75t_R   g4282( .A (y3198), .B (n4289), .Y (y1821) );
  AND3x1_ASAP7_75t_R   g4283( .A (n276), .B (x3), .C (x1), .Y (n4291) );
  OR3x1_ASAP7_75t_R    g4284( .A (n4291), .B (n81), .C (n10), .Y (y1822) );
  AO21x1_ASAP7_75t_R   g4285( .A1 (x4), .A2 (n58), .B (n2843), .Y (n4293) );
  OR3x1_ASAP7_75t_R    g4286( .A (n518), .B (n17), .C (n12), .Y (n4294) );
  INVx1_ASAP7_75t_R    g4287( .A (n4294), .Y (n4295) );
  AO21x1_ASAP7_75t_R   g4288( .A1 (n17), .A2 (n4293), .B (n4295), .Y (y1823) );
  AO21x1_ASAP7_75t_R   g4289( .A1 (n3474), .A2 (n1342), .B (n3055), .Y (y1824) );
  NOR2x1_ASAP7_75t_R   g4290( .A (n360), .B (n352), .Y (n4298) );
  INVx1_ASAP7_75t_R    g4291( .A (n4298), .Y (n4299) );
  AND3x1_ASAP7_75t_R   g4292( .A (n189), .B (y1894), .C (y3293), .Y (n4300) );
  AND2x2_ASAP7_75t_R   g4293( .A (n4299), .B (n4300), .Y (y1825) );
  AO21x1_ASAP7_75t_R   g4294( .A1 (n22), .A2 (x0), .B (n325), .Y (n4302) );
  NAND2x1_ASAP7_75t_R  g4295( .A (n353), .B (n4302), .Y (y1826) );
  AND2x2_ASAP7_75t_R   g4296( .A (n369), .B (n352), .Y (n4304) );
  AO21x1_ASAP7_75t_R   g4297( .A1 (x0), .A2 (x3), .B (n22), .Y (n4305) );
  OR3x1_ASAP7_75t_R    g4298( .A (y2196), .B (n368), .C (x4), .Y (n4306) );
  OA21x2_ASAP7_75t_R   g4299( .A1 (n4304), .A2 (n4305), .B (n4306), .Y (y1827) );
  NOR2x1_ASAP7_75t_R   g4300( .A (x3), .B (n473), .Y (n4308) );
  OR3x1_ASAP7_75t_R    g4301( .A (n4308), .B (n676), .C (n58), .Y (y1829) );
  AO32x1_ASAP7_75t_R   g4302( .A1 (n22), .A2 (n583), .A3 (n125), .B1 (x4), .B2 (n3327), .Y (y1830) );
  AO21x1_ASAP7_75t_R   g4303( .A1 (n29), .A2 (n77), .B (n529), .Y (y1831) );
  AO21x1_ASAP7_75t_R   g4304( .A1 (n90), .A2 (n22), .B (n537), .Y (n4312) );
  INVx1_ASAP7_75t_R    g4305( .A (n4312), .Y (n4313) );
  NAND2x1_ASAP7_75t_R  g4306( .A (y2079), .B (n3404), .Y (n4314) );
  OA21x2_ASAP7_75t_R   g4307( .A1 (n4313), .A2 (n4314), .B (n3712), .Y (y1832) );
  OA21x2_ASAP7_75t_R   g4308( .A1 (n4225), .A2 (n374), .B (y3377), .Y (y1833) );
  AO21x1_ASAP7_75t_R   g4309( .A1 (n360), .A2 (n290), .B (x2), .Y (n4317) );
  AND2x2_ASAP7_75t_R   g4310( .A (n4317), .B (n3029), .Y (y1834) );
  AO21x1_ASAP7_75t_R   g4311( .A1 (n596), .A2 (y2079), .B (n300), .Y (y1835) );
  AO21x1_ASAP7_75t_R   g4312( .A1 (n12), .A2 (n17), .B (y2466), .Y (n4320) );
  INVx1_ASAP7_75t_R    g4313( .A (n4320), .Y (n4321) );
  AO21x1_ASAP7_75t_R   g4314( .A1 (n4321), .A2 (n3119), .B (n344), .Y (y1836) );
  AO32x1_ASAP7_75t_R   g4315( .A1 (x0), .A2 (n22), .A3 (n319), .B1 (x4), .B2 (n3193), .Y (y1837) );
  NOR2x1_ASAP7_75t_R   g4316( .A (n589), .B (n1927), .Y (y1838) );
  OR3x1_ASAP7_75t_R    g4317( .A (n3027), .B (y2079), .C (n17), .Y (n4325) );
  AND2x2_ASAP7_75t_R   g4318( .A (n388), .B (n137), .Y (n4326) );
  NAND2x1_ASAP7_75t_R  g4319( .A (n4325), .B (n4326), .Y (y1839) );
  OA21x2_ASAP7_75t_R   g4320( .A1 (y1191), .A2 (n1454), .B (n1289), .Y (y1840) );
  OR3x1_ASAP7_75t_R    g4321( .A (n368), .B (x4), .C (x2), .Y (n4329) );
  AND2x2_ASAP7_75t_R   g4322( .A (n4329), .B (n3919), .Y (y1841) );
  OR3x1_ASAP7_75t_R    g4323( .A (y2022), .B (n22), .C (n43), .Y (n4331) );
  OA211x2_ASAP7_75t_R  g4324( .A1 (n3802), .A2 (x4), .B (n1782), .C (n4331), .Y (y1842) );
  AND3x1_ASAP7_75t_R   g4325( .A (n1586), .B (n762), .C (n86), .Y (y1843) );
  OA21x2_ASAP7_75t_R   g4326( .A1 (n628), .A2 (n300), .B (n3290), .Y (y1844) );
  AND3x1_ASAP7_75t_R   g4327( .A (n12), .B (n22), .C (x3), .Y (n4335) );
  INVx1_ASAP7_75t_R    g4328( .A (n4335), .Y (n4336) );
  AO32x1_ASAP7_75t_R   g4329( .A1 (y2079), .A2 (n4336), .A3 (n3620), .B1 (n22), .B2 (n3192), .Y (y1846) );
  OR3x1_ASAP7_75t_R    g4330( .A (n418), .B (x0), .C (x1), .Y (n4338) );
  AND3x1_ASAP7_75t_R   g4331( .A (n1717), .B (n4338), .C (y3293), .Y (y1847) );
  AND3x1_ASAP7_75t_R   g4332( .A (x2), .B (x4), .C (x5), .Y (n4340) );
  INVx1_ASAP7_75t_R    g4333( .A (n4340), .Y (n4341) );
  AND3x1_ASAP7_75t_R   g4334( .A (n4341), .B (n72), .C (n401), .Y (y1848) );
  AND3x1_ASAP7_75t_R   g4335( .A (n1110), .B (n3327), .C (n645), .Y (y1849) );
  AND2x2_ASAP7_75t_R   g4336( .A (n3380), .B (n219), .Y (y1850) );
  AND2x2_ASAP7_75t_R   g4337( .A (y195), .B (n1453), .Y (y1851) );
  AO21x1_ASAP7_75t_R   g4338( .A1 (n45), .A2 (n22), .B (y2079), .Y (y3527) );
  AND2x2_ASAP7_75t_R   g4339( .A (y3527), .B (n382), .Y (y1852) );
  AND2x2_ASAP7_75t_R   g4340( .A (n1970), .B (n3380), .Y (y1853) );
  AND3x1_ASAP7_75t_R   g4341( .A (n58), .B (n22), .C (n17), .Y (n4349) );
  AO21x1_ASAP7_75t_R   g4342( .A1 (n3291), .A2 (y2079), .B (n4349), .Y (y1854) );
  INVx1_ASAP7_75t_R    g4343( .A (n3160), .Y (n4351) );
  AO21x1_ASAP7_75t_R   g4344( .A1 (n4351), .A2 (n310), .B (n300), .Y (y1855) );
  OR3x1_ASAP7_75t_R    g4345( .A (y2466), .B (x3), .C (x0), .Y (n4353) );
  AND2x2_ASAP7_75t_R   g4346( .A (n4065), .B (n4353), .Y (y1856) );
  AND3x1_ASAP7_75t_R   g4347( .A (n152), .B (n153), .C (n1457), .Y (y1857) );
  AO21x1_ASAP7_75t_R   g4348( .A1 (n989), .A2 (n746), .B (n736), .Y (y1858) );
  AO21x1_ASAP7_75t_R   g4349( .A1 (n437), .A2 (x0), .B (y2079), .Y (n4357) );
  AND2x2_ASAP7_75t_R   g4350( .A (n906), .B (n4357), .Y (y1859) );
  AO21x1_ASAP7_75t_R   g4351( .A1 (n1093), .A2 (n22), .B (n1907), .Y (y1860) );
  NOR2x1_ASAP7_75t_R   g4352( .A (n12), .B (n368), .Y (n4360) );
  NOR2x1_ASAP7_75t_R   g4353( .A (n518), .B (n671), .Y (n4361) );
  OR3x1_ASAP7_75t_R    g4354( .A (n368), .B (n12), .C (x4), .Y (n4362) );
  OA21x2_ASAP7_75t_R   g4355( .A1 (n4360), .A2 (n4361), .B (n4362), .Y (y1861) );
  INVx1_ASAP7_75t_R    g4356( .A (n3977), .Y (y1862) );
  AND2x2_ASAP7_75t_R   g4357( .A (n917), .B (n968), .Y (y1863) );
  AND3x1_ASAP7_75t_R   g4358( .A (n15), .B (y2079), .C (x4), .Y (n4366) );
  AO32x1_ASAP7_75t_R   g4359( .A1 (n369), .A2 (n1265), .A3 (n370), .B1 (x3), .B2 (n4366), .Y (y1864) );
  AO21x1_ASAP7_75t_R   g4360( .A1 (n360), .A2 (n290), .B (n12), .Y (n4368) );
  NAND2x1_ASAP7_75t_R  g4361( .A (x5), .B (n4368), .Y (y1865) );
  OA21x2_ASAP7_75t_R   g4362( .A1 (n3477), .A2 (x5), .B (n367), .Y (y1866) );
  AO21x1_ASAP7_75t_R   g4363( .A1 (x2), .A2 (x3), .B (n22), .Y (n4371) );
  NAND2x1_ASAP7_75t_R  g4364( .A (y2079), .B (n4371), .Y (n4372) );
  AND3x1_ASAP7_75t_R   g4365( .A (x2), .B (x3), .C (x4), .Y (n4373) );
  INVx1_ASAP7_75t_R    g4366( .A (n4373), .Y (n4374) );
  AO21x1_ASAP7_75t_R   g4367( .A1 (x3), .A2 (x4), .B (n15), .Y (n4375) );
  NAND2x1_ASAP7_75t_R  g4368( .A (n4375), .B (n3762), .Y (n4376) );
  INVx1_ASAP7_75t_R    g4369( .A (n4376), .Y (n4377) );
  AO32x1_ASAP7_75t_R   g4370( .A1 (n1062), .A2 (n4372), .A3 (n4374), .B1 (y2079), .B2 (n4377), .Y (y1867) );
  OA21x2_ASAP7_75t_R   g4371( .A1 (n1477), .A2 (n267), .B (n2217), .Y (y1868) );
  AO21x1_ASAP7_75t_R   g4372( .A1 (n12), .A2 (n16), .B (n392), .Y (n4380) );
  NOR2x1_ASAP7_75t_R   g4373( .A (n468), .B (n4380), .Y (y1869) );
  OR3x1_ASAP7_75t_R    g4374( .A (n45), .B (x5), .C (x4), .Y (n4382) );
  AND2x2_ASAP7_75t_R   g4375( .A (n4151), .B (n4382), .Y (n4383) );
  AND3x1_ASAP7_75t_R   g4376( .A (n4383), .B (n1838), .C (n556), .Y (y1870) );
  NAND2x1_ASAP7_75t_R  g4377( .A (n12), .B (n1528), .Y (y1871) );
  OA22x2_ASAP7_75t_R   g4378( .A1 (y2079), .A2 (n3520), .B1 (n58), .B2 (n3521), .Y (y1872) );
  AO21x1_ASAP7_75t_R   g4379( .A1 (x0), .A2 (n544), .B (n1312), .Y (n4387) );
  AO21x1_ASAP7_75t_R   g4380( .A1 (x2), .A2 (n1305), .B (n4387), .Y (y1874) );
  INVx1_ASAP7_75t_R    g4381( .A (n501), .Y (n4389) );
  AO21x1_ASAP7_75t_R   g4382( .A1 (n4389), .A2 (x0), .B (n529), .Y (y1875) );
  AND3x1_ASAP7_75t_R   g4383( .A (n2217), .B (n2218), .C (n9), .Y (y1877) );
  OR3x1_ASAP7_75t_R    g4384( .A (n418), .B (x1), .C (x0), .Y (n4392) );
  AND3x1_ASAP7_75t_R   g4385( .A (n469), .B (n4392), .C (y3293), .Y (y1878) );
  AND3x1_ASAP7_75t_R   g4386( .A (n4037), .B (n1062), .C (y3293), .Y (y1879) );
  AO21x1_ASAP7_75t_R   g4387( .A1 (n17), .A2 (x5), .B (n325), .Y (n4395) );
  AND2x2_ASAP7_75t_R   g4388( .A (n4395), .B (n718), .Y (y1880) );
  AND3x1_ASAP7_75t_R   g4389( .A (y1702), .B (y3852), .C (n660), .Y (y1881) );
  AND2x2_ASAP7_75t_R   g4390( .A (n733), .B (n833), .Y (y1882) );
  AND2x2_ASAP7_75t_R   g4391( .A (n497), .B (n746), .Y (n4399) );
  AO21x1_ASAP7_75t_R   g4392( .A1 (y435), .A2 (n4399), .B (n2292), .Y (y1883) );
  AO21x1_ASAP7_75t_R   g4393( .A1 (n12), .A2 (n16), .B (n999), .Y (n4401) );
  AO21x1_ASAP7_75t_R   g4394( .A1 (y2079), .A2 (n4401), .B (n914), .Y (y1884) );
  AND3x1_ASAP7_75t_R   g4395( .A (n315), .B (y2079), .C (x3), .Y (n4403) );
  NOR2x1_ASAP7_75t_R   g4396( .A (n518), .B (n4403), .Y (y1885) );
  AND2x2_ASAP7_75t_R   g4397( .A (y2578), .B (x0), .Y (y1886) );
  AO32x1_ASAP7_75t_R   g4398( .A1 (y2079), .A2 (n4289), .A3 (n2645), .B1 (n22), .B2 (n3192), .Y (y1887) );
  AND3x1_ASAP7_75t_R   g4399( .A (n1853), .B (n451), .C (y1281), .Y (y1888) );
  AO21x1_ASAP7_75t_R   g4400( .A1 (n4037), .A2 (y3293), .B (n4038), .Y (y1889) );
  AND3x1_ASAP7_75t_R   g4401( .A (n455), .B (n137), .C (n72), .Y (n4409) );
  NAND2x1_ASAP7_75t_R  g4402( .A (n292), .B (n4409), .Y (y1890) );
  AND3x1_ASAP7_75t_R   g4403( .A (n401), .B (n583), .C (n3376), .Y (n4411) );
  INVx1_ASAP7_75t_R    g4404( .A (n4411), .Y (n4412) );
  AND2x2_ASAP7_75t_R   g4405( .A (n4412), .B (n3274), .Y (y1892) );
  AO21x1_ASAP7_75t_R   g4406( .A1 (n352), .A2 (n3085), .B (n3726), .Y (y1893) );
  AND3x1_ASAP7_75t_R   g4407( .A (n15), .B (x5), .C (x4), .Y (n4415) );
  INVx1_ASAP7_75t_R    g4408( .A (n4415), .Y (n4416) );
  AO21x1_ASAP7_75t_R   g4409( .A1 (y3293), .A2 (x2), .B (n4415), .Y (n4417) );
  AO32x1_ASAP7_75t_R   g4410( .A1 (n3780), .A2 (n4416), .A3 (n17), .B1 (x3), .B2 (n4417), .Y (y1895) );
  OR3x1_ASAP7_75t_R    g4411( .A (n211), .B (y2079), .C (x4), .Y (n4419) );
  INVx1_ASAP7_75t_R    g4412( .A (n4419), .Y (n4420) );
  AO21x1_ASAP7_75t_R   g4413( .A1 (n401), .A2 (n1269), .B (n4420), .Y (y1896) );
  OR3x1_ASAP7_75t_R    g4414( .A (n481), .B (y2196), .C (n15), .Y (n4422) );
  OR3x1_ASAP7_75t_R    g4415( .A (n58), .B (x2), .C (x1), .Y (n4423) );
  AND3x1_ASAP7_75t_R   g4416( .A (n4422), .B (n4423), .C (n144), .Y (n4424) );
  INVx1_ASAP7_75t_R    g4417( .A (n4424), .Y (y1897) );
  INVx1_ASAP7_75t_R    g4418( .A (n1815), .Y (n4426) );
  AO21x1_ASAP7_75t_R   g4419( .A1 (n228), .A2 (n1269), .B (n4426), .Y (y1898) );
  AO21x1_ASAP7_75t_R   g4420( .A1 (n262), .A2 (x3), .B (n81), .Y (y1899) );
  OR3x1_ASAP7_75t_R    g4421( .A (n856), .B (n12), .C (x1), .Y (n4429) );
  AND2x2_ASAP7_75t_R   g4422( .A (n4429), .B (n1424), .Y (y1900) );
  AND2x2_ASAP7_75t_R   g4423( .A (n72), .B (y2079), .Y (n4431) );
  AND3x1_ASAP7_75t_R   g4424( .A (n3469), .B (n3567), .C (n17), .Y (n4432) );
  INVx1_ASAP7_75t_R    g4425( .A (n4432), .Y (n4433) );
  OA21x2_ASAP7_75t_R   g4426( .A1 (n4431), .A2 (n3316), .B (n4433), .Y (y1901) );
  AO21x1_ASAP7_75t_R   g4427( .A1 (n337), .A2 (y2079), .B (x0), .Y (y3074) );
  AND2x2_ASAP7_75t_R   g4428( .A (y3074), .B (y3293), .Y (y1902) );
  AO21x1_ASAP7_75t_R   g4429( .A1 (n4116), .A2 (n22), .B (n3234), .Y (y1904) );
  AO21x1_ASAP7_75t_R   g4430( .A1 (y2079), .A2 (x2), .B (n3294), .Y (n4438) );
  AO21x1_ASAP7_75t_R   g4431( .A1 (n17), .A2 (x2), .B (n22), .Y (n4439) );
  AND2x2_ASAP7_75t_R   g4432( .A (n4438), .B (n4439), .Y (y1905) );
  NAND2x1_ASAP7_75t_R  g4433( .A (n406), .B (n3144), .Y (n4441) );
  AO21x1_ASAP7_75t_R   g4434( .A1 (n4441), .A2 (y1267), .B (y2466), .Y (y1906) );
  INVx1_ASAP7_75t_R    g4435( .A (n3338), .Y (n4443) );
  OR3x1_ASAP7_75t_R    g4436( .A (n4443), .B (n638), .C (x2), .Y (n4444) );
  AND2x2_ASAP7_75t_R   g4437( .A (n4444), .B (n4241), .Y (y1907) );
  AO21x1_ASAP7_75t_R   g4438( .A1 (n3979), .A2 (y2079), .B (n3085), .Y (y1908) );
  OA21x2_ASAP7_75t_R   g4439( .A1 (n3105), .A2 (n1319), .B (n556), .Y (y1909) );
  AND3x1_ASAP7_75t_R   g4440( .A (n58), .B (n17), .C (x4), .Y (n4448) );
  AO21x1_ASAP7_75t_R   g4441( .A1 (n2776), .A2 (n3148), .B (n4448), .Y (y1910) );
  OA21x2_ASAP7_75t_R   g4442( .A1 (n678), .A2 (x2), .B (n3919), .Y (y1911) );
  INVx1_ASAP7_75t_R    g4443( .A (n3193), .Y (n4451) );
  AOI22x1_ASAP7_75t_R  g4444( .A1 (n22), .A2 (n3193), .B1 (n4451), .B2 (n310), .Y (y1912) );
  AO21x1_ASAP7_75t_R   g4445( .A1 (x1), .A2 (n276), .B (n207), .Y (n4453) );
  AO32x1_ASAP7_75t_R   g4446( .A1 (n17), .A2 (n206), .A3 (n3955), .B1 (n145), .B2 (n4453), .Y (y1913) );
  AND3x1_ASAP7_75t_R   g4447( .A (n221), .B (y2079), .C (n15), .Y (n4455) );
  AO21x1_ASAP7_75t_R   g4448( .A1 (n232), .A2 (x2), .B (n4455), .Y (y1914) );
  AO21x1_ASAP7_75t_R   g4449( .A1 (n349), .A2 (x2), .B (n347), .Y (n4457) );
  AO21x1_ASAP7_75t_R   g4450( .A1 (n2979), .A2 (n4457), .B (n2982), .Y (y1915) );
  AND2x2_ASAP7_75t_R   g4451( .A (n3282), .B (y2079), .Y (n4459) );
  INVx1_ASAP7_75t_R    g4452( .A (n4070), .Y (n4460) );
  AO21x1_ASAP7_75t_R   g4453( .A1 (n4459), .A2 (n1572), .B (n4460), .Y (y1916) );
  AND3x1_ASAP7_75t_R   g4454( .A (n453), .B (y3852), .C (n466), .Y (y1917) );
  AO21x1_ASAP7_75t_R   g4455( .A1 (n576), .A2 (n1851), .B (x3), .Y (n4463) );
  AND2x2_ASAP7_75t_R   g4456( .A (n4463), .B (n3645), .Y (y1918) );
  AO21x1_ASAP7_75t_R   g4457( .A1 (n1062), .A2 (n3567), .B (n337), .Y (n4465) );
  NAND2x1_ASAP7_75t_R  g4458( .A (n4465), .B (n3584), .Y (y1919) );
  AO21x1_ASAP7_75t_R   g4459( .A1 (x3), .A2 (x2), .B (x5), .Y (n4467) );
  OA21x2_ASAP7_75t_R   g4460( .A1 (n3135), .A2 (n4243), .B (n4467), .Y (y1920) );
  OR3x1_ASAP7_75t_R    g4461( .A (n76), .B (x5), .C (x4), .Y (n4469) );
  NAND2x1_ASAP7_75t_R  g4462( .A (n4070), .B (n3794), .Y (y2739) );
  AND2x2_ASAP7_75t_R   g4463( .A (n4469), .B (y2739), .Y (y1921) );
  AO21x1_ASAP7_75t_R   g4464( .A1 (n129), .A2 (n58), .B (n1248), .Y (y1922) );
  AO21x1_ASAP7_75t_R   g4465( .A1 (n2504), .A2 (n1469), .B (n143), .Y (y1923) );
  AND3x1_ASAP7_75t_R   g4466( .A (n64), .B (n2158), .C (y2079), .Y (y1924) );
  AO21x1_ASAP7_75t_R   g4467( .A1 (n137), .A2 (n72), .B (n392), .Y (n4475) );
  INVx1_ASAP7_75t_R    g4468( .A (n4475), .Y (y1925) );
  AO21x1_ASAP7_75t_R   g4469( .A1 (n913), .A2 (n971), .B (n1184), .Y (y1926) );
  AO21x1_ASAP7_75t_R   g4470( .A1 (n12), .A2 (x5), .B (n403), .Y (n4478) );
  AND3x1_ASAP7_75t_R   g4471( .A (n378), .B (y3852), .C (n352), .Y (n4479) );
  AO21x1_ASAP7_75t_R   g4472( .A1 (y1702), .A2 (n4478), .B (n4479), .Y (y1927) );
  AO21x1_ASAP7_75t_R   g4473( .A1 (n559), .A2 (n1469), .B (n2169), .Y (y1928) );
  OR3x1_ASAP7_75t_R    g4474( .A (n337), .B (n15), .C (x5), .Y (n4482) );
  INVx1_ASAP7_75t_R    g4475( .A (n4482), .Y (n4483) );
  AO21x1_ASAP7_75t_R   g4476( .A1 (n22), .A2 (n3909), .B (n4483), .Y (y1929) );
  NOR2x1_ASAP7_75t_R   g4477( .A (n3118), .B (n3116), .Y (y1930) );
  INVx1_ASAP7_75t_R    g4478( .A (y3377), .Y (n4486) );
  AND3x1_ASAP7_75t_R   g4479( .A (n360), .B (n290), .C (n12), .Y (n4487) );
  NOR2x1_ASAP7_75t_R   g4480( .A (n4486), .B (n4487), .Y (y1931) );
  INVx1_ASAP7_75t_R    g4481( .A (n4401), .Y (n4489) );
  AND3x1_ASAP7_75t_R   g4482( .A (n968), .B (n219), .C (n419), .Y (n4490) );
  AO21x1_ASAP7_75t_R   g4483( .A1 (n1775), .A2 (n4489), .B (n4490), .Y (y1932) );
  OA21x2_ASAP7_75t_R   g4484( .A1 (n3963), .A2 (n22), .B (n3448), .Y (y1933) );
  AND2x2_ASAP7_75t_R   g4485( .A (y1635), .B (y1894), .Y (y1934) );
  INVx1_ASAP7_75t_R    g4486( .A (n3001), .Y (n4494) );
  AO21x1_ASAP7_75t_R   g4487( .A1 (n22), .A2 (x3), .B (n15), .Y (n4495) );
  AO21x1_ASAP7_75t_R   g4488( .A1 (n4494), .A2 (n4495), .B (n529), .Y (y1935) );
  AND2x2_ASAP7_75t_R   g4489( .A (n401), .B (n3469), .Y (n4497) );
  AO21x1_ASAP7_75t_R   g4490( .A1 (n4497), .A2 (y2079), .B (n3527), .Y (y1936) );
  AO21x1_ASAP7_75t_R   g4491( .A1 (n4497), .A2 (y2079), .B (n3847), .Y (y1937) );
  AO21x1_ASAP7_75t_R   g4492( .A1 (y2079), .A2 (n125), .B (n4349), .Y (y1938) );
  AO32x1_ASAP7_75t_R   g4493( .A1 (n17), .A2 (n2298), .A3 (n1490), .B1 (n185), .B2 (n259), .Y (y1939) );
  AO21x1_ASAP7_75t_R   g4494( .A1 (y2079), .A2 (x4), .B (n45), .Y (n4502) );
  AO21x1_ASAP7_75t_R   g4495( .A1 (n3568), .A2 (x5), .B (n4502), .Y (y3340) );
  NAND2x1_ASAP7_75t_R  g4496( .A (n15), .B (n641), .Y (n4504) );
  AND2x2_ASAP7_75t_R   g4497( .A (y3340), .B (n4504), .Y (y1940) );
  AO21x1_ASAP7_75t_R   g4498( .A1 (n1269), .A2 (n401), .B (n3847), .Y (y1941) );
  NAND2x1_ASAP7_75t_R  g4499( .A (x5), .B (n2992), .Y (n4507) );
  INVx1_ASAP7_75t_R    g4500( .A (n641), .Y (n4508) );
  AND2x2_ASAP7_75t_R   g4501( .A (n4507), .B (n4508), .Y (y1942) );
  AND3x1_ASAP7_75t_R   g4502( .A (n2116), .B (n2117), .C (y2079), .Y (y1943) );
  AO21x1_ASAP7_75t_R   g4503( .A1 (n1062), .A2 (n660), .B (n3183), .Y (y1944) );
  OA222x2_ASAP7_75t_R  g4504( .A1 (n3182), .A2 (n3585), .B1 (n22), .B2 (y2079), .C1 (n3181), .C2 (n3584), .Y (y1945) );
  OA21x2_ASAP7_75t_R   g4505( .A1 (n29), .A2 (n4401), .B (y3852), .Y (y1946) );
  AND3x1_ASAP7_75t_R   g4506( .A (n22), .B (n17), .C (x5), .Y (n4514) );
  AO21x1_ASAP7_75t_R   g4507( .A1 (y2079), .A2 (n348), .B (n4514), .Y (n4515) );
  AND2x2_ASAP7_75t_R   g4508( .A (n4515), .B (n330), .Y (y1947) );
  AND3x1_ASAP7_75t_R   g4509( .A (n2211), .B (n219), .C (n64), .Y (y1948) );
  INVx1_ASAP7_75t_R    g4510( .A (n4375), .Y (n4518) );
  OR3x1_ASAP7_75t_R    g4511( .A (n4518), .B (y2079), .C (n3333), .Y (n4519) );
  NAND2x1_ASAP7_75t_R  g4512( .A (x2), .B (n641), .Y (n4520) );
  AND2x2_ASAP7_75t_R   g4513( .A (n4519), .B (n4520), .Y (y1949) );
  AO21x1_ASAP7_75t_R   g4514( .A1 (n67), .A2 (n703), .B (n2347), .Y (y1950) );
  NAND2x1_ASAP7_75t_R  g4515( .A (n316), .B (n310), .Y (n4523) );
  AND2x2_ASAP7_75t_R   g4516( .A (n4523), .B (n3290), .Y (y1951) );
  AND2x2_ASAP7_75t_R   g4517( .A (n770), .B (n707), .Y (y1952) );
  AO21x1_ASAP7_75t_R   g4518( .A1 (n17), .A2 (x4), .B (x5), .Y (n4526) );
  INVx1_ASAP7_75t_R    g4519( .A (n4526), .Y (n4527) );
  AO21x1_ASAP7_75t_R   g4520( .A1 (x4), .A2 (x5), .B (x2), .Y (n4528) );
  NOR2x1_ASAP7_75t_R   g4521( .A (x3), .B (n4528), .Y (n4529) );
  AO21x1_ASAP7_75t_R   g4522( .A1 (n4527), .A2 (x2), .B (n4529), .Y (y1953) );
  AO21x1_ASAP7_75t_R   g4523( .A1 (y2079), .A2 (n511), .B (n300), .Y (y1954) );
  NAND2x1_ASAP7_75t_R  g4524( .A (n316), .B (n3567), .Y (n4532) );
  AO21x1_ASAP7_75t_R   g4525( .A1 (n45), .A2 (n455), .B (n4532), .Y (y1955) );
  OA21x2_ASAP7_75t_R   g4526( .A1 (n1269), .A2 (n1457), .B (n770), .Y (y1956) );
  AND3x1_ASAP7_75t_R   g4527( .A (n17), .B (x4), .C (x2), .Y (n4535) );
  INVx1_ASAP7_75t_R    g4528( .A (n4535), .Y (n4536) );
  AO32x1_ASAP7_75t_R   g4529( .A1 (y2079), .A2 (n4536), .A3 (n3377), .B1 (n337), .B2 (n1646), .Y (y1957) );
  NAND2x1_ASAP7_75t_R  g4530( .A (n1980), .B (n976), .Y (y1958) );
  AO21x1_ASAP7_75t_R   g4531( .A1 (n173), .A2 (n1646), .B (y2163), .Y (y1959) );
  NAND2x1_ASAP7_75t_R  g4532( .A (y2079), .B (n334), .Y (n4540) );
  INVx1_ASAP7_75t_R    g4533( .A (n4540), .Y (n4541) );
  AO21x1_ASAP7_75t_R   g4534( .A1 (n22), .A2 (n3191), .B (n4541), .Y (y1960) );
  AO21x1_ASAP7_75t_R   g4535( .A1 (n90), .A2 (n750), .B (n839), .Y (n4543) );
  AND2x2_ASAP7_75t_R   g4536( .A (n4543), .B (n244), .Y (y1961) );
  AO21x1_ASAP7_75t_R   g4537( .A1 (n84), .A2 (n125), .B (n22), .Y (n4545) );
  AND3x1_ASAP7_75t_R   g4538( .A (n3977), .B (n4545), .C (n3327), .Y (y1962) );
  NAND2x1_ASAP7_75t_R  g4539( .A (n18), .B (n1527), .Y (y1963) );
  OR3x1_ASAP7_75t_R    g4540( .A (n529), .B (n29), .C (n15), .Y (n4548) );
  OA21x2_ASAP7_75t_R   g4541( .A1 (x2), .A2 (n1277), .B (n4548), .Y (y1964) );
  AND2x2_ASAP7_75t_R   g4542( .A (n3469), .B (n3567), .Y (n4550) );
  INVx1_ASAP7_75t_R    g4543( .A (n4550), .Y (n4551) );
  AND2x2_ASAP7_75t_R   g4544( .A (n3001), .B (n2998), .Y (n4552) );
  AO21x1_ASAP7_75t_R   g4545( .A1 (n4551), .A2 (n17), .B (n4552), .Y (y1965) );
  AND3x1_ASAP7_75t_R   g4546( .A (n189), .B (n369), .C (x4), .Y (n4554) );
  AO21x1_ASAP7_75t_R   g4547( .A1 (n125), .A2 (n29), .B (n4554), .Y (y1966) );
  AND2x2_ASAP7_75t_R   g4548( .A (y201), .B (n52), .Y (y1967) );
  NAND2x1_ASAP7_75t_R  g4549( .A (n4232), .B (n740), .Y (y1968) );
  AO21x1_ASAP7_75t_R   g4550( .A1 (n52), .A2 (n58), .B (n716), .Y (y1969) );
  AO21x1_ASAP7_75t_R   g4551( .A1 (n299), .A2 (n310), .B (n672), .Y (n4559) );
  AND2x2_ASAP7_75t_R   g4552( .A (y3198), .B (n4559), .Y (y1970) );
  AO21x1_ASAP7_75t_R   g4553( .A1 (n28), .A2 (x3), .B (n3237), .Y (n4561) );
  INVx1_ASAP7_75t_R    g4554( .A (n4561), .Y (n4562) );
  AO21x1_ASAP7_75t_R   g4555( .A1 (n3237), .A2 (n4443), .B (n4562), .Y (y1971) );
  NOR2x1_ASAP7_75t_R   g4556( .A (n22), .B (n756), .Y (n4564) );
  AO21x1_ASAP7_75t_R   g4557( .A1 (n660), .A2 (n1062), .B (n4564), .Y (y1972) );
  AND3x1_ASAP7_75t_R   g4558( .A (n217), .B (n406), .C (n632), .Y (y1973) );
  AO21x1_ASAP7_75t_R   g4559( .A1 (y2079), .A2 (x4), .B (n3279), .Y (n4567) );
  AO21x1_ASAP7_75t_R   g4560( .A1 (n45), .A2 (n28), .B (n4567), .Y (y1974) );
  INVx1_ASAP7_75t_R    g4561( .A (n3909), .Y (n4569) );
  AND3x1_ASAP7_75t_R   g4562( .A (n4569), .B (n388), .C (n360), .Y (n4570) );
  INVx1_ASAP7_75t_R    g4563( .A (n4570), .Y (n4571) );
  AND2x2_ASAP7_75t_R   g4564( .A (x5), .B (x3), .Y (n4572) );
  AO21x1_ASAP7_75t_R   g4565( .A1 (n4572), .A2 (x4), .B (x2), .Y (n4573) );
  AND2x2_ASAP7_75t_R   g4566( .A (n4571), .B (n4573), .Y (y1975) );
  INVx1_ASAP7_75t_R    g4567( .A (n3794), .Y (n4575) );
  AND3x1_ASAP7_75t_R   g4568( .A (n17), .B (n15), .C (x5), .Y (n4576) );
  OA21x2_ASAP7_75t_R   g4569( .A1 (n4575), .A2 (n4576), .B (n2998), .Y (y1976) );
  AND3x1_ASAP7_75t_R   g4570( .A (n1265), .B (n3023), .C (n290), .Y (y1977) );
  AND3x1_ASAP7_75t_R   g4571( .A (y1393), .B (n906), .C (n899), .Y (y1978) );
  NOR2x1_ASAP7_75t_R   g4572( .A (x5), .B (n176), .Y (y1979) );
  AO21x1_ASAP7_75t_R   g4573( .A1 (x1), .A2 (n537), .B (n512), .Y (n4581) );
  OR3x1_ASAP7_75t_R    g4574( .A (n4581), .B (n29), .C (n529), .Y (y1980) );
  AO21x1_ASAP7_75t_R   g4575( .A1 (x4), .A2 (n12), .B (n319), .Y (n4583) );
  INVx1_ASAP7_75t_R    g4576( .A (n4583), .Y (n4584) );
  OR3x1_ASAP7_75t_R    g4577( .A (n4584), .B (n3129), .C (n914), .Y (y1981) );
  AND3x1_ASAP7_75t_R   g4578( .A (n22), .B (y2079), .C (x3), .Y (n4586) );
  NOR2x1_ASAP7_75t_R   g4579( .A (n4586), .B (n3301), .Y (n4587) );
  NAND2x1_ASAP7_75t_R  g4580( .A (n15), .B (n4099), .Y (n4588) );
  INVx1_ASAP7_75t_R    g4581( .A (n4588), .Y (n4589) );
  AO21x1_ASAP7_75t_R   g4582( .A1 (n4587), .A2 (x2), .B (n4589), .Y (y1982) );
  AO21x1_ASAP7_75t_R   g4583( .A1 (x2), .A2 (n403), .B (n3316), .Y (n4591) );
  AND2x2_ASAP7_75t_R   g4584( .A (n4591), .B (n2971), .Y (y1983) );
  AO32x1_ASAP7_75t_R   g4585( .A1 (n3524), .A2 (x5), .A3 (n3000), .B1 (n3567), .B2 (n3585), .Y (y1984) );
  OR3x1_ASAP7_75t_R    g4586( .A (n418), .B (n15), .C (n17), .Y (n4594) );
  AO21x1_ASAP7_75t_R   g4587( .A1 (n17), .A2 (n15), .B (n392), .Y (n4595) );
  INVx1_ASAP7_75t_R    g4588( .A (n4595), .Y (n4596) );
  AND2x2_ASAP7_75t_R   g4589( .A (n4594), .B (n4596), .Y (y1985) );
  AO21x1_ASAP7_75t_R   g4590( .A1 (x2), .A2 (x4), .B (n17), .Y (n4598) );
  AND3x1_ASAP7_75t_R   g4591( .A (n757), .B (n290), .C (n4598), .Y (y1986) );
  AO21x1_ASAP7_75t_R   g4592( .A1 (n40), .A2 (n228), .B (n2099), .Y (y1987) );
  AO21x1_ASAP7_75t_R   g4593( .A1 (n12), .A2 (x1), .B (x3), .Y (n4601) );
  INVx1_ASAP7_75t_R    g4594( .A (n4601), .Y (n4602) );
  AO21x1_ASAP7_75t_R   g4595( .A1 (n4602), .A2 (n1469), .B (n2581), .Y (y1988) );
  AND3x1_ASAP7_75t_R   g4596( .A (n1269), .B (n360), .C (n290), .Y (n4604) );
  AO21x1_ASAP7_75t_R   g4597( .A1 (n337), .A2 (n1646), .B (n4604), .Y (y1989) );
  NAND2x1_ASAP7_75t_R  g4598( .A (x2), .B (n3800), .Y (n4606) );
  AO21x1_ASAP7_75t_R   g4599( .A1 (n3800), .A2 (x2), .B (n164), .Y (n4607) );
  AO32x1_ASAP7_75t_R   g4600( .A1 (n72), .A2 (n4606), .A3 (y435), .B1 (n221), .B2 (n4607), .Y (n4608) );
  INVx1_ASAP7_75t_R    g4601( .A (n4608), .Y (y1990) );
  AO21x1_ASAP7_75t_R   g4602( .A1 (n1646), .A2 (n377), .B (n4137), .Y (y1991) );
  AO21x1_ASAP7_75t_R   g4603( .A1 (y2079), .A2 (x2), .B (n403), .Y (n4611) );
  AO21x1_ASAP7_75t_R   g4604( .A1 (n97), .A2 (n740), .B (n337), .Y (n4612) );
  AOI22x1_ASAP7_75t_R  g4605( .A1 (n378), .A2 (n1646), .B1 (n4611), .B2 (n4612), .Y (y1992) );
  AO21x1_ASAP7_75t_R   g4606( .A1 (n22), .A2 (x1), .B (n967), .Y (n4614) );
  AND2x2_ASAP7_75t_R   g4607( .A (n4614), .B (y2079), .Y (n4615) );
  NOR2x1_ASAP7_75t_R   g4608( .A (n3748), .B (n4615), .Y (y1993) );
  NOR2x1_ASAP7_75t_R   g4609( .A (n3859), .B (n3989), .Y (y1994) );
  INVx1_ASAP7_75t_R    g4610( .A (n3598), .Y (n4618) );
  AO21x1_ASAP7_75t_R   g4611( .A1 (x5), .A2 (x4), .B (x3), .Y (n4619) );
  AND3x1_ASAP7_75t_R   g4612( .A (n4618), .B (n4619), .C (n3148), .Y (y1995) );
  INVx1_ASAP7_75t_R    g4613( .A (n3905), .Y (n4621) );
  AND2x2_ASAP7_75t_R   g4614( .A (n4109), .B (n3944), .Y (y2015) );
  OA21x2_ASAP7_75t_R   g4615( .A1 (x3), .A2 (n4621), .B (y2015), .Y (y1996) );
  AO21x1_ASAP7_75t_R   g4616( .A1 (n219), .A2 (n90), .B (y1891), .Y (y1998) );
  INVx1_ASAP7_75t_R    g4617( .A (n994), .Y (n4625) );
  AND3x1_ASAP7_75t_R   g4618( .A (y3852), .B (n994), .C (x4), .Y (n4626) );
  AO21x1_ASAP7_75t_R   g4619( .A1 (n492), .A2 (n4625), .B (n4626), .Y (n4627) );
  AO21x1_ASAP7_75t_R   g4620( .A1 (x0), .A2 (x1), .B (n4627), .Y (y1999) );
  AND2x2_ASAP7_75t_R   g4621( .A (n3924), .B (n1971), .Y (y2000) );
  OA21x2_ASAP7_75t_R   g4622( .A1 (x2), .A2 (n337), .B (n3285), .Y (y2001) );
  NOR2x1_ASAP7_75t_R   g4623( .A (x3), .B (n3011), .Y (n4631) );
  INVx1_ASAP7_75t_R    g4624( .A (n4631), .Y (n4632) );
  OR3x1_ASAP7_75t_R    g4625( .A (n45), .B (n22), .C (y2079), .Y (n4633) );
  AND2x2_ASAP7_75t_R   g4626( .A (n4632), .B (n4633), .Y (y2002) );
  AO21x1_ASAP7_75t_R   g4627( .A1 (n12), .A2 (x4), .B (n17), .Y (n4635) );
  NAND2x1_ASAP7_75t_R  g4628( .A (n3267), .B (n4635), .Y (n4636) );
  OA21x2_ASAP7_75t_R   g4629( .A1 (n4636), .A2 (x5), .B (y3198), .Y (y2003) );
  OR3x1_ASAP7_75t_R    g4630( .A (x3), .B (x2), .C (x5), .Y (n4638) );
  AO32x1_ASAP7_75t_R   g4631( .A1 (n22), .A2 (n217), .A3 (n319), .B1 (n4638), .B2 (n4243), .Y (y2004) );
  NAND2x1_ASAP7_75t_R  g4632( .A (n388), .B (n3567), .Y (n4640) );
  AO32x1_ASAP7_75t_R   g4633( .A1 (n388), .A2 (n3272), .A3 (n3567), .B1 (n672), .B2 (n4640), .Y (y2005) );
  AND2x2_ASAP7_75t_R   g4634( .A (y1903), .B (n3797), .Y (y2006) );
  OR3x1_ASAP7_75t_R    g4635( .A (n325), .B (n15), .C (x5), .Y (n4643) );
  INVx1_ASAP7_75t_R    g4636( .A (n4643), .Y (n4644) );
  AO21x1_ASAP7_75t_R   g4637( .A1 (y2740), .A2 (n15), .B (n4644), .Y (y2007) );
  AND2x2_ASAP7_75t_R   g4638( .A (y1393), .B (n1385), .Y (y2008) );
  AO21x1_ASAP7_75t_R   g4639( .A1 (n137), .A2 (n72), .B (n22), .Y (n4647) );
  INVx1_ASAP7_75t_R    g4640( .A (n4647), .Y (n4648) );
  NOR2x1_ASAP7_75t_R   g4641( .A (n3992), .B (n4648), .Y (n4649) );
  NOR2x1_ASAP7_75t_R   g4642( .A (n4486), .B (n4649), .Y (y2009) );
  OR3x1_ASAP7_75t_R    g4643( .A (n211), .B (x5), .C (x4), .Y (n4651) );
  AO21x1_ASAP7_75t_R   g4644( .A1 (n15), .A2 (y2079), .B (n4250), .Y (y2882) );
  AND2x2_ASAP7_75t_R   g4645( .A (n4651), .B (y2882), .Y (y2010) );
  AO21x1_ASAP7_75t_R   g4646( .A1 (n16), .A2 (x4), .B (n58), .Y (n4654) );
  OA21x2_ASAP7_75t_R   g4647( .A1 (n1078), .A2 (n4654), .B (n919), .Y (y2011) );
  INVx1_ASAP7_75t_R    g4648( .A (n2559), .Y (n4656) );
  AND3x1_ASAP7_75t_R   g4649( .A (n3955), .B (y9), .C (n17), .Y (n4657) );
  AO21x1_ASAP7_75t_R   g4650( .A1 (n4656), .A2 (x3), .B (n4657), .Y (y2012) );
  OR3x1_ASAP7_75t_R    g4651( .A (n3073), .B (n2718), .C (n29), .Y (y2013) );
  AO21x1_ASAP7_75t_R   g4652( .A1 (n22), .A2 (n4467), .B (n4648), .Y (n4660) );
  AND2x2_ASAP7_75t_R   g4653( .A (n4660), .B (n2971), .Y (y2014) );
  OR3x1_ASAP7_75t_R    g4654( .A (n58), .B (n17), .C (x4), .Y (n4662) );
  OA21x2_ASAP7_75t_R   g4655( .A1 (n3112), .A2 (n22), .B (n4662), .Y (y2017) );
  AO32x1_ASAP7_75t_R   g4656( .A1 (y3293), .A2 (n1062), .A3 (n391), .B1 (n3584), .B2 (n3182), .Y (y2018) );
  AO21x1_ASAP7_75t_R   g4657( .A1 (x4), .A2 (x2), .B (n17), .Y (n4665) );
  AO21x1_ASAP7_75t_R   g4658( .A1 (n22), .A2 (n15), .B (x3), .Y (n4666) );
  NAND2x1_ASAP7_75t_R  g4659( .A (n4665), .B (n4666), .Y (n4667) );
  AO21x1_ASAP7_75t_R   g4660( .A1 (n81), .A2 (n22), .B (y2079), .Y (n4668) );
  OA21x2_ASAP7_75t_R   g4661( .A1 (n4667), .A2 (x5), .B (n4668), .Y (y2019) );
  INVx1_ASAP7_75t_R    g4662( .A (n478), .Y (n4670) );
  AO21x1_ASAP7_75t_R   g4663( .A1 (n4670), .A2 (n23), .B (n529), .Y (y2020) );
  AND2x2_ASAP7_75t_R   g4664( .A (n348), .B (y3852), .Y (n4672) );
  AND2x2_ASAP7_75t_R   g4665( .A (n3647), .B (n4672), .Y (y2021) );
  AO21x1_ASAP7_75t_R   g4666( .A1 (n2999), .A2 (n17), .B (y2079), .Y (n4674) );
  AND3x1_ASAP7_75t_R   g4667( .A (n3625), .B (n4674), .C (n660), .Y (y2023) );
  AND3x1_ASAP7_75t_R   g4668( .A (n217), .B (n2117), .C (y9), .Y (y3963) );
  AO21x1_ASAP7_75t_R   g4669( .A1 (n16), .A2 (n812), .B (y3963), .Y (y2024) );
  INVx1_ASAP7_75t_R    g4670( .A (n389), .Y (n4678) );
  AO21x1_ASAP7_75t_R   g4671( .A1 (n17), .A2 (x0), .B (y2466), .Y (n4679) );
  AND2x2_ASAP7_75t_R   g4672( .A (n4678), .B (n4679), .Y (y2025) );
  INVx1_ASAP7_75t_R    g4673( .A (n2051), .Y (n4681) );
  AND2x2_ASAP7_75t_R   g4674( .A (n4681), .B (y3527), .Y (y2026) );
  AO21x1_ASAP7_75t_R   g4675( .A1 (n12), .A2 (n16), .B (n243), .Y (n4683) );
  INVx1_ASAP7_75t_R    g4676( .A (n4683), .Y (n4684) );
  OA21x2_ASAP7_75t_R   g4677( .A1 (n4684), .A2 (n276), .B (n2729), .Y (y2027) );
  AOI21x1_ASAP7_75t_R  g4678( .A1 (n3825), .A2 (n3824), .B (n392), .Y (y2028) );
  AND2x2_ASAP7_75t_R   g4679( .A (n968), .B (n604), .Y (y2029) );
  AO21x1_ASAP7_75t_R   g4680( .A1 (n17), .A2 (x4), .B (n12), .Y (n4688) );
  AO21x1_ASAP7_75t_R   g4681( .A1 (n421), .A2 (n22), .B (x0), .Y (n4689) );
  OA21x2_ASAP7_75t_R   g4682( .A1 (n366), .A2 (n4688), .B (n4689), .Y (y2030) );
  AND2x2_ASAP7_75t_R   g4683( .A (n3023), .B (n4439), .Y (y2031) );
  OA21x2_ASAP7_75t_R   g4684( .A1 (x4), .A2 (n1210), .B (n496), .Y (y2032) );
  INVx1_ASAP7_75t_R    g4685( .A (n4529), .Y (n4693) );
  OR3x1_ASAP7_75t_R    g4686( .A (n45), .B (y2079), .C (n22), .Y (y3397) );
  AO21x1_ASAP7_75t_R   g4687( .A1 (x2), .A2 (x5), .B (x4), .Y (n4695) );
  AND3x1_ASAP7_75t_R   g4688( .A (n4693), .B (y3397), .C (n4695), .Y (y2033) );
  AND2x2_ASAP7_75t_R   g4689( .A (n4302), .B (n3579), .Y (y2035) );
  AO32x1_ASAP7_75t_R   g4690( .A1 (n316), .A2 (n3028), .A3 (n3618), .B1 (x2), .B2 (n628), .Y (y2036) );
  AND2x2_ASAP7_75t_R   g4691( .A (n129), .B (n244), .Y (n4699) );
  OA21x2_ASAP7_75t_R   g4692( .A1 (n4699), .A2 (n2914), .B (n2360), .Y (y2037) );
  NOR2x1_ASAP7_75t_R   g4693( .A (x5), .B (n4487), .Y (y2038) );
  AO21x1_ASAP7_75t_R   g4694( .A1 (n15), .A2 (x5), .B (n231), .Y (n4702) );
  INVx1_ASAP7_75t_R    g4695( .A (n4702), .Y (n4703) );
  OA33x2_ASAP7_75t_R   g4696( .A1 (n231), .A2 (n1646), .A3 (y772), .B1 (n746), .B2 (n4703), .B3 (n993), .Y (y2039) );
  AO21x1_ASAP7_75t_R   g4697( .A1 (x4), .A2 (n3294), .B (n3592), .Y (y2040) );
  OR3x1_ASAP7_75t_R    g4698( .A (n2544), .B (n2546), .C (n109), .Y (y2041) );
  AND2x2_ASAP7_75t_R   g4699( .A (n3579), .B (n3267), .Y (y2042) );
  AO21x1_ASAP7_75t_R   g4700( .A1 (x3), .A2 (x5), .B (n22), .Y (n4708) );
  AND2x2_ASAP7_75t_R   g4701( .A (n369), .B (n740), .Y (n4709) );
  OAI22x1_ASAP7_75t_R  g4702( .A1 (n4708), .A2 (n4180), .B1 (n4709), .B2 (x4), .Y (y2043) );
  NAND2x1_ASAP7_75t_R  g4703( .A (n292), .B (n3181), .Y (y2044) );
  AND3x1_ASAP7_75t_R   g4704( .A (n3660), .B (n382), .C (y2079), .Y (y3633) );
  AO21x1_ASAP7_75t_R   g4705( .A1 (n22), .A2 (n421), .B (y3633), .Y (y2045) );
  NAND2x1_ASAP7_75t_R  g4706( .A (n3040), .B (n652), .Y (n4714) );
  AND2x2_ASAP7_75t_R   g4707( .A (n4714), .B (y3377), .Y (y2046) );
  AO21x1_ASAP7_75t_R   g4708( .A1 (n125), .A2 (n474), .B (n4554), .Y (y2047) );
  AO32x1_ASAP7_75t_R   g4709( .A1 (n84), .A2 (n352), .A3 (n22), .B1 (n2645), .B2 (y2079), .Y (y2048) );
  AND2x2_ASAP7_75t_R   g4710( .A (n1870), .B (n1247), .Y (y2049) );
  AND3x1_ASAP7_75t_R   g4711( .A (n221), .B (y2079), .C (n22), .Y (n4719) );
  INVx1_ASAP7_75t_R    g4712( .A (n4719), .Y (n4720) );
  NAND2x1_ASAP7_75t_R  g4713( .A (x5), .B (n1707), .Y (y2632) );
  AND2x2_ASAP7_75t_R   g4714( .A (n4720), .B (y2632), .Y (y2050) );
  AO21x1_ASAP7_75t_R   g4715( .A1 (n12), .A2 (y2079), .B (n368), .Y (n4723) );
  AO21x1_ASAP7_75t_R   g4716( .A1 (n22), .A2 (n4723), .B (n4554), .Y (y2051) );
  AND2x2_ASAP7_75t_R   g4717( .A (n496), .B (n4670), .Y (y2052) );
  NAND2x1_ASAP7_75t_R  g4718( .A (n22), .B (n4200), .Y (n4726) );
  INVx1_ASAP7_75t_R    g4719( .A (n4576), .Y (n4727) );
  AND3x1_ASAP7_75t_R   g4720( .A (n4726), .B (n3794), .C (n4727), .Y (n4728) );
  INVx1_ASAP7_75t_R    g4721( .A (n4728), .Y (y2053) );
  NOR2x1_ASAP7_75t_R   g4722( .A (n2600), .B (n4486), .Y (y2054) );
  AND3x1_ASAP7_75t_R   g4723( .A (n12), .B (x1), .C (x4), .Y (n4731) );
  INVx1_ASAP7_75t_R    g4724( .A (n4731), .Y (n4732) );
  AO21x1_ASAP7_75t_R   g4725( .A1 (n4732), .A2 (n972), .B (n3572), .Y (y2055) );
  AO21x1_ASAP7_75t_R   g4726( .A1 (n290), .A2 (n360), .B (n15), .Y (n4734) );
  AND3x1_ASAP7_75t_R   g4727( .A (n3927), .B (n4734), .C (n556), .Y (y2056) );
  AO21x1_ASAP7_75t_R   g4728( .A1 (y2079), .A2 (x4), .B (n337), .Y (n4736) );
  AO21x1_ASAP7_75t_R   g4729( .A1 (x0), .A2 (x5), .B (x3), .Y (n4737) );
  AND2x2_ASAP7_75t_R   g4730( .A (n4736), .B (n4737), .Y (y2057) );
  INVx1_ASAP7_75t_R    g4731( .A (n809), .Y (n4739) );
  AO21x1_ASAP7_75t_R   g4732( .A1 (n4739), .A2 (n12), .B (y863), .Y (n4740) );
  AO21x1_ASAP7_75t_R   g4733( .A1 (n4740), .A2 (n217), .B (n222), .Y (y2058) );
  AO21x1_ASAP7_75t_R   g4734( .A1 (y2079), .A2 (n401), .B (n3751), .Y (y2059) );
  AO21x1_ASAP7_75t_R   g4735( .A1 (n4219), .A2 (n1191), .B (n344), .Y (y2060) );
  AND2x2_ASAP7_75t_R   g4736( .A (n3469), .B (n3023), .Y (y2061) );
  NAND2x1_ASAP7_75t_R  g4737( .A (n1106), .B (y3852), .Y (n4745) );
  XOR2x2_ASAP7_75t_R   g4738( .A (n4745), .B (n916), .Y (y2062) );
  AO21x1_ASAP7_75t_R   g4739( .A1 (n1163), .A2 (n3327), .B (n3009), .Y (y2063) );
  NAND2x1_ASAP7_75t_R  g4740( .A (x0), .B (n464), .Y (n4748) );
  OA21x2_ASAP7_75t_R   g4741( .A1 (x0), .A2 (n552), .B (n4748), .Y (y2064) );
  OA21x2_ASAP7_75t_R   g4742( .A1 (n3603), .A2 (y2079), .B (n3924), .Y (y2065) );
  AO21x1_ASAP7_75t_R   g4743( .A1 (n22), .A2 (n17), .B (n76), .Y (n4751) );
  AND2x2_ASAP7_75t_R   g4744( .A (n4751), .B (n3237), .Y (y2066) );
  AO21x1_ASAP7_75t_R   g4745( .A1 (n22), .A2 (y2079), .B (n15), .Y (n4753) );
  INVx1_ASAP7_75t_R    g4746( .A (n4753), .Y (n4754) );
  OR3x1_ASAP7_75t_R    g4747( .A (n529), .B (n29), .C (n17), .Y (n4755) );
  AO32x1_ASAP7_75t_R   g4748( .A1 (x3), .A2 (n396), .A3 (n4753), .B1 (n4754), .B2 (n4755), .Y (y2067) );
  NAND2x1_ASAP7_75t_R  g4749( .A (x2), .B (n2576), .Y (n4757) );
  AO21x1_ASAP7_75t_R   g4750( .A1 (n13), .A2 (x0), .B (n17), .Y (n4758) );
  AND2x2_ASAP7_75t_R   g4751( .A (n4757), .B (n4758), .Y (y2069) );
  AO21x1_ASAP7_75t_R   g4752( .A1 (y2079), .A2 (n125), .B (n3085), .Y (y2070) );
  OA21x2_ASAP7_75t_R   g4753( .A1 (n3568), .A2 (n45), .B (n3029), .Y (y2071) );
  AO21x1_ASAP7_75t_R   g4754( .A1 (y2079), .A2 (n22), .B (y570), .Y (y2072) );
  AO21x1_ASAP7_75t_R   g4755( .A1 (n90), .A2 (n17), .B (n120), .Y (n4763) );
  AO21x1_ASAP7_75t_R   g4756( .A1 (n16), .A2 (x0), .B (x3), .Y (n4764) );
  INVx1_ASAP7_75t_R    g4757( .A (n4764), .Y (n4765) );
  NAND2x1_ASAP7_75t_R  g4758( .A (n15), .B (n4765), .Y (n4766) );
  AOI21x1_ASAP7_75t_R  g4759( .A1 (n4763), .A2 (n4766), .B (n1208), .Y (y2073) );
  AND3x1_ASAP7_75t_R   g4760( .A (n401), .B (n1265), .C (n3376), .Y (n4768) );
  NOR2x1_ASAP7_75t_R   g4761( .A (n3624), .B (n4768), .Y (y2074) );
  NOR2x1_ASAP7_75t_R   g4762( .A (n386), .B (n3434), .Y (y2075) );
  INVx1_ASAP7_75t_R    g4763( .A (n4024), .Y (n4771) );
  AND2x2_ASAP7_75t_R   g4764( .A (n3446), .B (n77), .Y (y2274) );
  OA21x2_ASAP7_75t_R   g4765( .A1 (n4771), .A2 (y2274), .B (n3987), .Y (y2076) );
  AO21x1_ASAP7_75t_R   g4766( .A1 (n413), .A2 (y2079), .B (n3189), .Y (y2077) );
  AO21x1_ASAP7_75t_R   g4767( .A1 (n17), .A2 (n15), .B (y2466), .Y (n4775) );
  AND2x2_ASAP7_75t_R   g4768( .A (n3678), .B (n4775), .Y (y2078) );
  AO32x1_ASAP7_75t_R   g4769( .A1 (n17), .A2 (n3013), .A3 (n3011), .B1 (n22), .B2 (y2079), .Y (n4777) );
  AO21x1_ASAP7_75t_R   g4770( .A1 (n164), .A2 (y3293), .B (n4777), .Y (y2080) );
  AND3x1_ASAP7_75t_R   g4771( .A (n3797), .B (y1281), .C (n3979), .Y (y2081) );
  NAND2x1_ASAP7_75t_R  g4772( .A (n45), .B (n388), .Y (n4780) );
  INVx1_ASAP7_75t_R    g4773( .A (n4780), .Y (n4781) );
  OR3x1_ASAP7_75t_R    g4774( .A (n4781), .B (n3867), .C (n3568), .Y (y2082) );
  AND2x2_ASAP7_75t_R   g4775( .A (y0), .B (y2079), .Y (y2083) );
  AND3x1_ASAP7_75t_R   g4776( .A (n173), .B (n174), .C (x3), .Y (n4784) );
  AO21x1_ASAP7_75t_R   g4777( .A1 (x0), .A2 (n103), .B (n4784), .Y (y2084) );
  AO21x1_ASAP7_75t_R   g4778( .A1 (x3), .A2 (n22), .B (n3327), .Y (y2085) );
  AND2x2_ASAP7_75t_R   g4779( .A (n369), .B (n4305), .Y (y2086) );
  AND3x1_ASAP7_75t_R   g4780( .A (n15), .B (y2079), .C (x3), .Y (n4788) );
  INVx1_ASAP7_75t_R    g4781( .A (n4788), .Y (n4789) );
  AND3x1_ASAP7_75t_R   g4782( .A (n3943), .B (n4789), .C (n556), .Y (y2087) );
  AO21x1_ASAP7_75t_R   g4783( .A1 (n757), .A2 (n4136), .B (n4137), .Y (y2088) );
  AND3x1_ASAP7_75t_R   g4784( .A (n45), .B (n22), .C (x5), .Y (n4792) );
  AO21x1_ASAP7_75t_R   g4785( .A1 (x4), .A2 (n3611), .B (n4792), .Y (y2089) );
  NOR2x1_ASAP7_75t_R   g4786( .A (x5), .B (n950), .Y (y2090) );
  AND2x2_ASAP7_75t_R   g4787( .A (n2524), .B (n707), .Y (n4795) );
  OA21x2_ASAP7_75t_R   g4788( .A1 (n16), .A2 (n2508), .B (n4795), .Y (y2091) );
  AO32x1_ASAP7_75t_R   g4789( .A1 (n1265), .A2 (n3944), .A3 (x3), .B1 (x4), .B2 (n4709), .Y (y2092) );
  AND2x2_ASAP7_75t_R   g4790( .A (y3397), .B (n3024), .Y (y2094) );
  AO21x1_ASAP7_75t_R   g4791( .A1 (n63), .A2 (n363), .B (n754), .Y (y2095) );
  AO21x1_ASAP7_75t_R   g4792( .A1 (n2470), .A2 (x1), .B (n1644), .Y (y2096) );
  AO21x1_ASAP7_75t_R   g4793( .A1 (n352), .A2 (n337), .B (n3234), .Y (y2097) );
  AND3x1_ASAP7_75t_R   g4794( .A (y3198), .B (n3797), .C (n660), .Y (y2098) );
  AND2x2_ASAP7_75t_R   g4795( .A (y2740), .B (n583), .Y (y2099) );
  AND2x2_ASAP7_75t_R   g4796( .A (n3804), .B (n4070), .Y (n4804) );
  AND3x1_ASAP7_75t_R   g4797( .A (n4804), .B (n77), .C (y2079), .Y (y2100) );
  AND3x1_ASAP7_75t_R   g4798( .A (n1370), .B (n1196), .C (n219), .Y (y2101) );
  AO21x1_ASAP7_75t_R   g4799( .A1 (n628), .A2 (n1851), .B (n638), .Y (y2102) );
  NOR2x1_ASAP7_75t_R   g4800( .A (x5), .B (n1150), .Y (n4808) );
  AO21x1_ASAP7_75t_R   g4801( .A1 (n3365), .A2 (n970), .B (n4808), .Y (y2103) );
  AO21x1_ASAP7_75t_R   g4802( .A1 (n427), .A2 (n22), .B (n529), .Y (y2104) );
  NAND2x1_ASAP7_75t_R  g4803( .A (y2079), .B (y25), .Y (n4811) );
  INVx1_ASAP7_75t_R    g4804( .A (n4811), .Y (y2105) );
  AO21x1_ASAP7_75t_R   g4805( .A1 (n1209), .A2 (n15), .B (n2169), .Y (y2106) );
  OA21x2_ASAP7_75t_R   g4806( .A1 (n993), .A2 (n1851), .B (n3380), .Y (y2107) );
  INVx1_ASAP7_75t_R    g4807( .A (n2104), .Y (n4815) );
  AND2x2_ASAP7_75t_R   g4808( .A (y3852), .B (n290), .Y (n4816) );
  NAND2x1_ASAP7_75t_R  g4809( .A (x3), .B (n718), .Y (n4817) );
  AND2x2_ASAP7_75t_R   g4810( .A (n4816), .B (n4817), .Y (n4818) );
  NOR2x1_ASAP7_75t_R   g4811( .A (n4815), .B (n4818), .Y (y2108) );
  AND3x1_ASAP7_75t_R   g4812( .A (x2), .B (x4), .C (x3), .Y (n4820) );
  INVx1_ASAP7_75t_R    g4813( .A (n4820), .Y (n4821) );
  AO21x1_ASAP7_75t_R   g4814( .A1 (n4821), .A2 (n348), .B (y2079), .Y (n4822) );
  OA211x2_ASAP7_75t_R  g4815( .A1 (n285), .A2 (n4820), .B (n4822), .C (n2980), .Y (y2109) );
  AO21x1_ASAP7_75t_R   g4816( .A1 (y3293), .A2 (x3), .B (n1277), .Y (n4824) );
  AND3x1_ASAP7_75t_R   g4817( .A (n4824), .B (n419), .C (x0), .Y (y2110) );
  OA21x2_ASAP7_75t_R   g4818( .A1 (n1032), .A2 (n337), .B (y3852), .Y (y2111) );
  AND2x2_ASAP7_75t_R   g4819( .A (n652), .B (y2079), .Y (y2112) );
  AO21x1_ASAP7_75t_R   g4820( .A1 (n2542), .A2 (n1209), .B (n1208), .Y (n4828) );
  NAND2x1_ASAP7_75t_R  g4821( .A (n388), .B (n4828), .Y (y2113) );
  OR3x1_ASAP7_75t_R    g4822( .A (n518), .B (n17), .C (n15), .Y (n4830) );
  INVx1_ASAP7_75t_R    g4823( .A (n4830), .Y (n4831) );
  AO21x1_ASAP7_75t_R   g4824( .A1 (n28), .A2 (n45), .B (n4831), .Y (y2114) );
  OR3x1_ASAP7_75t_R    g4825( .A (n3384), .B (n3386), .C (x5), .Y (n4833) );
  AND2x2_ASAP7_75t_R   g4826( .A (n4833), .B (y2135), .Y (y2115) );
  INVx1_ASAP7_75t_R    g4827( .A (n4349), .Y (n4835) );
  OA21x2_ASAP7_75t_R   g4828( .A1 (n3005), .A2 (n22), .B (n4835), .Y (y2116) );
  AO21x1_ASAP7_75t_R   g4829( .A1 (n1775), .A2 (x3), .B (n4349), .Y (y2117) );
  AO21x1_ASAP7_75t_R   g4830( .A1 (n378), .A2 (x0), .B (y2740), .Y (y2118) );
  AND2x2_ASAP7_75t_R   g4831( .A (n3968), .B (n556), .Y (y2119) );
  AO21x1_ASAP7_75t_R   g4832( .A1 (n137), .A2 (y2079), .B (n756), .Y (n4840) );
  AND2x2_ASAP7_75t_R   g4833( .A (n3278), .B (x4), .Y (n4841) );
  AO21x1_ASAP7_75t_R   g4834( .A1 (n22), .A2 (n4840), .B (n4841), .Y (y2120) );
  AND3x1_ASAP7_75t_R   g4835( .A (n17), .B (x5), .C (x2), .Y (n4843) );
  AO21x1_ASAP7_75t_R   g4836( .A1 (n15), .A2 (x3), .B (x4), .Y (n4844) );
  OA21x2_ASAP7_75t_R   g4837( .A1 (n4843), .A2 (n4844), .B (n3907), .Y (y2121) );
  AO21x1_ASAP7_75t_R   g4838( .A1 (n669), .A2 (x0), .B (n344), .Y (y2122) );
  INVx1_ASAP7_75t_R    g4839( .A (n2847), .Y (n4847) );
  AO21x1_ASAP7_75t_R   g4840( .A1 (n4847), .A2 (n144), .B (n2169), .Y (y2123) );
  AO21x1_ASAP7_75t_R   g4841( .A1 (y2079), .A2 (x3), .B (n3294), .Y (n4849) );
  AND2x2_ASAP7_75t_R   g4842( .A (n4022), .B (n22), .Y (n4850) );
  XOR2x2_ASAP7_75t_R   g4843( .A (n4849), .B (n4850), .Y (y2124) );
  OA21x2_ASAP7_75t_R   g4844( .A1 (n1128), .A2 (n604), .B (n1102), .Y (y2125) );
  AO21x1_ASAP7_75t_R   g4845( .A1 (y3852), .A2 (n22), .B (n781), .Y (n4853) );
  AND3x1_ASAP7_75t_R   g4846( .A (n1211), .B (n4853), .C (n556), .Y (y2126) );
  AO21x1_ASAP7_75t_R   g4847( .A1 (n90), .A2 (x2), .B (n826), .Y (n4855) );
  INVx1_ASAP7_75t_R    g4848( .A (n4855), .Y (n4856) );
  AO21x1_ASAP7_75t_R   g4849( .A1 (n4856), .A2 (n17), .B (n2581), .Y (y2127) );
  AND3x1_ASAP7_75t_R   g4850( .A (y3198), .B (n3128), .C (n3797), .Y (y2128) );
  AO21x1_ASAP7_75t_R   g4851( .A1 (y2079), .A2 (n299), .B (n989), .Y (y2129) );
  NOR2x1_ASAP7_75t_R   g4852( .A (x5), .B (n374), .Y (y2130) );
  NOR2x1_ASAP7_75t_R   g4853( .A (n16), .B (n2738), .Y (n4861) );
  AO21x1_ASAP7_75t_R   g4854( .A1 (n797), .A2 (n120), .B (n4861), .Y (y2131) );
  AND2x2_ASAP7_75t_R   g4855( .A (n3057), .B (n1720), .Y (y2132) );
  AO21x1_ASAP7_75t_R   g4856( .A1 (x4), .A2 (n58), .B (y2466), .Y (n4864) );
  AO21x1_ASAP7_75t_R   g4857( .A1 (n622), .A2 (n4864), .B (n399), .Y (y2133) );
  AO21x1_ASAP7_75t_R   g4858( .A1 (y9), .A2 (y2466), .B (n143), .Y (y2134) );
  AO21x1_ASAP7_75t_R   g4859( .A1 (y2079), .A2 (n360), .B (n914), .Y (y2136) );
  INVx1_ASAP7_75t_R    g4860( .A (n4232), .Y (n4868) );
  OA21x2_ASAP7_75t_R   g4861( .A1 (n286), .A2 (n4868), .B (n382), .Y (y2137) );
  AND3x1_ASAP7_75t_R   g4862( .A (n451), .B (n3327), .C (n290), .Y (y2138) );
  AND2x2_ASAP7_75t_R   g4863( .A (n2366), .B (n2182), .Y (y2139) );
  AO21x1_ASAP7_75t_R   g4864( .A1 (y3377), .A2 (n724), .B (n4225), .Y (y2140) );
  AO21x1_ASAP7_75t_R   g4865( .A1 (n15), .A2 (n1245), .B (n2527), .Y (y2141) );
  NAND2x1_ASAP7_75t_R  g4866( .A (n415), .B (n3520), .Y (n4874) );
  AND2x2_ASAP7_75t_R   g4867( .A (n4874), .B (y2079), .Y (y2142) );
  INVx1_ASAP7_75t_R    g4868( .A (n3896), .Y (n4876) );
  AO21x1_ASAP7_75t_R   g4869( .A1 (n15), .A2 (x3), .B (n3027), .Y (n4877) );
  NOR2x1_ASAP7_75t_R   g4870( .A (n406), .B (n4877), .Y (n4878) );
  AO21x1_ASAP7_75t_R   g4871( .A1 (y2079), .A2 (n4876), .B (n4878), .Y (y2143) );
  OA21x2_ASAP7_75t_R   g4872( .A1 (n4015), .A2 (y2196), .B (n645), .Y (y2145) );
  AO21x1_ASAP7_75t_R   g4873( .A1 (n4426), .A2 (n22), .B (n529), .Y (y2146) );
  NAND2x1_ASAP7_75t_R  g4874( .A (n4070), .B (n3804), .Y (n4882) );
  AO21x1_ASAP7_75t_R   g4875( .A1 (n3804), .A2 (n4070), .B (y2079), .Y (y3386) );
  OA21x2_ASAP7_75t_R   g4876( .A1 (n4882), .A2 (x5), .B (y3386), .Y (y2148) );
  AO21x1_ASAP7_75t_R   g4877( .A1 (n17), .A2 (n583), .B (n425), .Y (n4885) );
  AO32x1_ASAP7_75t_R   g4878( .A1 (n1431), .A2 (n1434), .A3 (n529), .B1 (n22), .B2 (n4885), .Y (y2149) );
  AO21x1_ASAP7_75t_R   g4879( .A1 (n382), .A2 (x0), .B (n2051), .Y (y3556) );
  AND2x2_ASAP7_75t_R   g4880( .A (y3556), .B (n3212), .Y (y2150) );
  AO21x1_ASAP7_75t_R   g4881( .A1 (n143), .A2 (x2), .B (n17), .Y (n4889) );
  AND2x2_ASAP7_75t_R   g4882( .A (n2814), .B (n4889), .Y (y2151) );
  AND2x2_ASAP7_75t_R   g4883( .A (n497), .B (n219), .Y (n4891) );
  OR3x1_ASAP7_75t_R    g4884( .A (n495), .B (n978), .C (x2), .Y (n4892) );
  OA21x2_ASAP7_75t_R   g4885( .A1 (n4891), .A2 (n15), .B (n4892), .Y (y2152) );
  AO21x1_ASAP7_75t_R   g4886( .A1 (x5), .A2 (n1150), .B (n1078), .Y (y2153) );
  AND3x1_ASAP7_75t_R   g4887( .A (n401), .B (n1265), .C (n3143), .Y (n4895) );
  AND2x2_ASAP7_75t_R   g4888( .A (n4895), .B (n4241), .Y (y2154) );
  OA21x2_ASAP7_75t_R   g4889( .A1 (n3085), .A2 (n3978), .B (n3327), .Y (y2156) );
  AO21x1_ASAP7_75t_R   g4890( .A1 (n495), .A2 (n22), .B (x0), .Y (n4898) );
  AND2x2_ASAP7_75t_R   g4891( .A (n600), .B (n4898), .Y (y2157) );
  AO21x1_ASAP7_75t_R   g4892( .A1 (n1191), .A2 (n1247), .B (n495), .Y (y2158) );
  AND3x1_ASAP7_75t_R   g4893( .A (n3028), .B (n3377), .C (y2079), .Y (y2159) );
  AND3x1_ASAP7_75t_R   g4894( .A (n3446), .B (n3448), .C (n2998), .Y (y2160) );
  AO21x1_ASAP7_75t_R   g4895( .A1 (y2079), .A2 (x3), .B (n22), .Y (n4903) );
  NAND2x1_ASAP7_75t_R  g4896( .A (n22), .B (n3285), .Y (n4904) );
  OA21x2_ASAP7_75t_R   g4897( .A1 (n3294), .A2 (n4903), .B (n4904), .Y (y2161) );
  AND2x2_ASAP7_75t_R   g4898( .A (y2740), .B (x0), .Y (y2162) );
  AO21x1_ASAP7_75t_R   g4899( .A1 (x5), .A2 (n22), .B (n125), .Y (n4907) );
  INVx1_ASAP7_75t_R    g4900( .A (n4907), .Y (n4908) );
  OR3x1_ASAP7_75t_R    g4901( .A (n399), .B (n4908), .C (n315), .Y (y2164) );
  AND3x1_ASAP7_75t_R   g4902( .A (n72), .B (n137), .C (n22), .Y (n4910) );
  INVx1_ASAP7_75t_R    g4903( .A (n4910), .Y (n4911) );
  AND2x2_ASAP7_75t_R   g4904( .A (n4911), .B (n3946), .Y (y2165) );
  NAND2x1_ASAP7_75t_R  g4905( .A (n312), .B (n310), .Y (y2166) );
  AO21x1_ASAP7_75t_R   g4906( .A1 (n72), .A2 (n137), .B (n22), .Y (n4914) );
  INVx1_ASAP7_75t_R    g4907( .A (n4914), .Y (n4915) );
  AO21x1_ASAP7_75t_R   g4908( .A1 (y2079), .A2 (x2), .B (x3), .Y (n4916) );
  INVx1_ASAP7_75t_R    g4909( .A (n4916), .Y (n4917) );
  OA21x2_ASAP7_75t_R   g4910( .A1 (n4917), .A2 (n3611), .B (n22), .Y (n4918) );
  AO21x1_ASAP7_75t_R   g4911( .A1 (n4915), .A2 (y2079), .B (n4918), .Y (y2167) );
  INVx1_ASAP7_75t_R    g4912( .A (n1319), .Y (n4920) );
  NAND2x1_ASAP7_75t_R  g4913( .A (x0), .B (n3443), .Y (n4921) );
  INVx1_ASAP7_75t_R    g4914( .A (n4921), .Y (n4922) );
  AO21x1_ASAP7_75t_R   g4915( .A1 (y3852), .A2 (n4920), .B (n4922), .Y (y2168) );
  AO21x1_ASAP7_75t_R   g4916( .A1 (n3469), .A2 (n3567), .B (x3), .Y (n4924) );
  INVx1_ASAP7_75t_R    g4917( .A (n4924), .Y (n4925) );
  AO21x1_ASAP7_75t_R   g4918( .A1 (n3029), .A2 (x3), .B (n4925), .Y (n4926) );
  AND2x2_ASAP7_75t_R   g4919( .A (n4926), .B (n1265), .Y (y2169) );
  AO21x1_ASAP7_75t_R   g4920( .A1 (n413), .A2 (n348), .B (n363), .Y (y2170) );
  AO21x1_ASAP7_75t_R   g4921( .A1 (n4754), .A2 (n366), .B (n45), .Y (y2171) );
  AND3x1_ASAP7_75t_R   g4922( .A (n2542), .B (n299), .C (y2079), .Y (y2172) );
  INVx1_ASAP7_75t_R    g4923( .A (y1702), .Y (n4931) );
  INVx1_ASAP7_75t_R    g4924( .A (n1997), .Y (n4932) );
  AO21x1_ASAP7_75t_R   g4925( .A1 (n299), .A2 (y2079), .B (n4932), .Y (n4933) );
  OA21x2_ASAP7_75t_R   g4926( .A1 (n4931), .A2 (n3376), .B (n4933), .Y (y2173) );
  OR3x1_ASAP7_75t_R    g4927( .A (n227), .B (x5), .C (x4), .Y (n4935) );
  AND3x1_ASAP7_75t_R   g4928( .A (n2986), .B (y2813), .C (n4935), .Y (y2174) );
  AO21x1_ASAP7_75t_R   g4929( .A1 (n12), .A2 (x1), .B (n15), .Y (n4937) );
  NAND2x1_ASAP7_75t_R  g4930( .A (n2038), .B (n4937), .Y (n4938) );
  AND2x2_ASAP7_75t_R   g4931( .A (n4938), .B (n1510), .Y (y2175) );
  NAND2x1_ASAP7_75t_R  g4932( .A (n139), .B (n388), .Y (n4940) );
  AND3x1_ASAP7_75t_R   g4933( .A (n4940), .B (n369), .C (n572), .Y (y2176) );
  NAND2x1_ASAP7_75t_R  g4934( .A (n3083), .B (n3567), .Y (n4942) );
  OA21x2_ASAP7_75t_R   g4935( .A1 (n4942), .A2 (n1158), .B (n3943), .Y (y2177) );
  AND3x1_ASAP7_75t_R   g4936( .A (n90), .B (n219), .C (n620), .Y (y2178) );
  AND2x2_ASAP7_75t_R   g4937( .A (n64), .B (y3852), .Y (n4945) );
  AND2x2_ASAP7_75t_R   g4938( .A (n2623), .B (n4945), .Y (y2179) );
  AO21x1_ASAP7_75t_R   g4939( .A1 (n3990), .A2 (y2079), .B (n3135), .Y (y2180) );
  INVx1_ASAP7_75t_R    g4940( .A (n2572), .Y (n4948) );
  AND3x1_ASAP7_75t_R   g4941( .A (n4948), .B (n4014), .C (n22), .Y (n4949) );
  AO21x1_ASAP7_75t_R   g4942( .A1 (x5), .A2 (n12), .B (n290), .Y (n4950) );
  INVx1_ASAP7_75t_R    g4943( .A (n4950), .Y (n4951) );
  OR3x1_ASAP7_75t_R    g4944( .A (n4949), .B (n4951), .C (y2196), .Y (y2181) );
  OR3x1_ASAP7_75t_R    g4945( .A (n403), .B (n15), .C (x5), .Y (n4953) );
  INVx1_ASAP7_75t_R    g4946( .A (n4953), .Y (n4954) );
  NOR2x1_ASAP7_75t_R   g4947( .A (n4954), .B (n3761), .Y (y2182) );
  AO331x2_ASAP7_75t_R  g4948( .A1 (x2), .A2 (n388), .A3 (n3338), .B1 (n15), .B2 (n401), .B3 (n3565), .C (n3443), .Y (y2183) );
  AO21x1_ASAP7_75t_R   g4949( .A1 (y2079), .A2 (n436), .B (n914), .Y (n4957) );
  AND2x2_ASAP7_75t_R   g4950( .A (n4957), .B (n1354), .Y (y2184) );
  AO21x1_ASAP7_75t_R   g4951( .A1 (y2079), .A2 (n17), .B (n22), .Y (n4959) );
  AO21x1_ASAP7_75t_R   g4952( .A1 (x5), .A2 (x3), .B (x2), .Y (n4960) );
  INVx1_ASAP7_75t_R    g4953( .A (n4960), .Y (n4961) );
  NAND2x1_ASAP7_75t_R  g4954( .A (n4959), .B (n4961), .Y (n4962) );
  AND3x1_ASAP7_75t_R   g4955( .A (n4962), .B (n3019), .C (n336), .Y (y2185) );
  AND3x1_ASAP7_75t_R   g4956( .A (n77), .B (n3804), .C (x5), .Y (n4964) );
  AO21x1_ASAP7_75t_R   g4957( .A1 (n1572), .A2 (n4459), .B (n4964), .Y (y2186) );
  AND3x1_ASAP7_75t_R   g4958( .A (y3198), .B (n3797), .C (n661), .Y (y2187) );
  AO21x1_ASAP7_75t_R   g4959( .A1 (n645), .A2 (n3327), .B (n3085), .Y (y2188) );
  NAND2x1_ASAP7_75t_R  g4960( .A (n4907), .B (n398), .Y (y2189) );
  AND2x2_ASAP7_75t_R   g4961( .A (y3758), .B (n218), .Y (y2771) );
  AO21x1_ASAP7_75t_R   g4962( .A1 (n4775), .A2 (n3860), .B (y2771), .Y (y2190) );
  AND3x1_ASAP7_75t_R   g4963( .A (n2141), .B (n2150), .C (n3091), .Y (y2191) );
  AO21x1_ASAP7_75t_R   g4964( .A1 (n17), .A2 (x4), .B (n15), .Y (n4972) );
  AO32x1_ASAP7_75t_R   g4965( .A1 (n740), .A2 (n4536), .A3 (n4598), .B1 (n4972), .B2 (n366), .Y (n4973) );
  INVx1_ASAP7_75t_R    g4966( .A (n4973), .Y (y2192) );
  AO21x1_ASAP7_75t_R   g4967( .A1 (y2079), .A2 (x3), .B (n4349), .Y (y2193) );
  AO21x1_ASAP7_75t_R   g4968( .A1 (x0), .A2 (x3), .B (n16), .Y (n4976) );
  AO21x1_ASAP7_75t_R   g4969( .A1 (n1296), .A2 (n4976), .B (n15), .Y (n4977) );
  AND3x1_ASAP7_75t_R   g4970( .A (n15), .B (x1), .C (x3), .Y (n4978) );
  INVx1_ASAP7_75t_R    g4971( .A (n4978), .Y (n4979) );
  AND2x2_ASAP7_75t_R   g4972( .A (n4977), .B (n4979), .Y (y2194) );
  NOR2x1_ASAP7_75t_R   g4973( .A (n15), .B (n368), .Y (n4981) );
  AO21x1_ASAP7_75t_R   g4974( .A1 (n15), .A2 (n368), .B (n4981), .Y (n4982) );
  NOR2x1_ASAP7_75t_R   g4975( .A (n22), .B (n4982), .Y (n4983) );
  NOR2x1_ASAP7_75t_R   g4976( .A (n4420), .B (n4983), .Y (y2195) );
  AO21x1_ASAP7_75t_R   g4977( .A1 (n22), .A2 (n3828), .B (n1269), .Y (y2197) );
  AO21x1_ASAP7_75t_R   g4978( .A1 (n4304), .A2 (n22), .B (n3234), .Y (y2198) );
  NAND2x1_ASAP7_75t_R  g4979( .A (n16), .B (n2060), .Y (n4987) );
  AND2x2_ASAP7_75t_R   g4980( .A (n4987), .B (n1455), .Y (y2199) );
  AND3x1_ASAP7_75t_R   g4981( .A (n1863), .B (y1281), .C (n1853), .Y (y2200) );
  OR3x1_ASAP7_75t_R    g4982( .A (n392), .B (n17), .C (n15), .Y (n4990) );
  INVx1_ASAP7_75t_R    g4983( .A (n4990), .Y (n4991) );
  AO21x1_ASAP7_75t_R   g4984( .A1 (n419), .A2 (n45), .B (n4991), .Y (y2201) );
  AND2x2_ASAP7_75t_R   g4985( .A (y232), .B (y2079), .Y (y2202) );
  AO21x1_ASAP7_75t_R   g4986( .A1 (y1656), .A2 (n2596), .B (n3974), .Y (y2203) );
  AO21x1_ASAP7_75t_R   g4987( .A1 (n3777), .A2 (x2), .B (n529), .Y (n4995) );
  AO21x1_ASAP7_75t_R   g4988( .A1 (n15), .A2 (n17), .B (n4995), .Y (y2204) );
  AO21x1_ASAP7_75t_R   g4989( .A1 (n84), .A2 (n29), .B (n3005), .Y (y2205) );
  INVx1_ASAP7_75t_R    g4990( .A (n1510), .Y (n4998) );
  NOR2x1_ASAP7_75t_R   g4991( .A (n4998), .B (n65), .Y (y2206) );
  NAND2x1_ASAP7_75t_R  g4992( .A (x5), .B (n4465), .Y (y3084) );
  AO21x1_ASAP7_75t_R   g4993( .A1 (x2), .A2 (x4), .B (x5), .Y (n5001) );
  AND2x2_ASAP7_75t_R   g4994( .A (y3084), .B (n5001), .Y (y2207) );
  AO21x1_ASAP7_75t_R   g4995( .A1 (y2079), .A2 (x0), .B (n139), .Y (n5003) );
  INVx1_ASAP7_75t_R    g4996( .A (n5003), .Y (n5004) );
  AO21x1_ASAP7_75t_R   g4997( .A1 (n5004), .A2 (n660), .B (n529), .Y (y2208) );
  NAND2x1_ASAP7_75t_R  g4998( .A (n3072), .B (n356), .Y (y2209) );
  INVx1_ASAP7_75t_R    g4999( .A (n4638), .Y (n5007) );
  AO21x1_ASAP7_75t_R   g5000( .A1 (n1572), .A2 (n455), .B (n3860), .Y (n5008) );
  AO21x1_ASAP7_75t_R   g5001( .A1 (n5007), .A2 (n22), .B (n5008), .Y (n5009) );
  INVx1_ASAP7_75t_R    g5002( .A (n5009), .Y (y2210) );
  AO21x1_ASAP7_75t_R   g5003( .A1 (n16), .A2 (n1646), .B (y1207), .Y (y2211) );
  NOR2x1_ASAP7_75t_R   g5004( .A (x5), .B (n3732), .Y (n5012) );
  AO32x1_ASAP7_75t_R   g5005( .A1 (n22), .A2 (y435), .A3 (n1242), .B1 (n228), .B2 (n5012), .Y (y2212) );
  OR3x1_ASAP7_75t_R    g5006( .A (n3637), .B (x5), .C (x3), .Y (n5014) );
  AND2x2_ASAP7_75t_R   g5007( .A (n5014), .B (n406), .Y (y2213) );
  AND3x1_ASAP7_75t_R   g5008( .A (n388), .B (n137), .C (n72), .Y (n5016) );
  INVx1_ASAP7_75t_R    g5009( .A (n3548), .Y (n5017) );
  NOR2x1_ASAP7_75t_R   g5010( .A (n5017), .B (n5016), .Y (y2815) );
  AO21x1_ASAP7_75t_R   g5011( .A1 (n5016), .A2 (n5017), .B (y2815), .Y (y2214) );
  AO32x1_ASAP7_75t_R   g5012( .A1 (n348), .A2 (n4129), .A3 (n757), .B1 (n17), .B2 (n3279), .Y (y2215) );
  AND2x2_ASAP7_75t_R   g5013( .A (y2134), .B (n556), .Y (y2216) );
  AND3x1_ASAP7_75t_R   g5014( .A (n241), .B (n17), .C (n16), .Y (n5022) );
  AO21x1_ASAP7_75t_R   g5015( .A1 (n1572), .A2 (n143), .B (n5022), .Y (y2217) );
  OA21x2_ASAP7_75t_R   g5016( .A1 (n421), .A2 (n4844), .B (n3907), .Y (y2218) );
  AND2x2_ASAP7_75t_R   g5017( .A (y2393), .B (y2079), .Y (y2221) );
  OR3x1_ASAP7_75t_R    g5018( .A (n271), .B (n262), .C (n227), .Y (y3802) );
  AND2x2_ASAP7_75t_R   g5019( .A (y3802), .B (y2079), .Y (y2222) );
  AO21x1_ASAP7_75t_R   g5020( .A1 (n90), .A2 (n219), .B (n1269), .Y (y2223) );
  AND2x2_ASAP7_75t_R   g5021( .A (n3977), .B (y1438), .Y (y2224) );
  AO21x1_ASAP7_75t_R   g5022( .A1 (n17), .A2 (y2079), .B (x2), .Y (n5030) );
  AO32x1_ASAP7_75t_R   g5023( .A1 (x4), .A2 (n672), .A3 (n3023), .B1 (n22), .B2 (n5030), .Y (y2225) );
  NAND2x1_ASAP7_75t_R  g5024( .A (x3), .B (n1391), .Y (n5032) );
  AND2x2_ASAP7_75t_R   g5025( .A (n5032), .B (n173), .Y (n5033) );
  NAND2x1_ASAP7_75t_R  g5026( .A (x2), .B (n184), .Y (n5034) );
  INVx1_ASAP7_75t_R    g5027( .A (n5034), .Y (n5035) );
  AOI21x1_ASAP7_75t_R  g5028( .A1 (n187), .A2 (n5033), .B (n5035), .Y (y2226) );
  INVx1_ASAP7_75t_R    g5029( .A (n4937), .Y (n5037) );
  OA21x2_ASAP7_75t_R   g5030( .A1 (n5037), .A2 (n145), .B (n1656), .Y (y2227) );
  NOR2x1_ASAP7_75t_R   g5031( .A (n3327), .B (n3072), .Y (n5039) );
  AND2x2_ASAP7_75t_R   g5032( .A (n3327), .B (n3072), .Y (n5040) );
  OR3x1_ASAP7_75t_R    g5033( .A (n5039), .B (n5040), .C (y2196), .Y (y2228) );
  AND3x1_ASAP7_75t_R   g5034( .A (y2632), .B (n1240), .C (n4935), .Y (y2229) );
  AO21x1_ASAP7_75t_R   g5035( .A1 (x3), .A2 (n3819), .B (n3899), .Y (y2230) );
  AO21x1_ASAP7_75t_R   g5036( .A1 (n1528), .A2 (x0), .B (n787), .Y (y2231) );
  AO21x1_ASAP7_75t_R   g5037( .A1 (n2971), .A2 (n4467), .B (n3316), .Y (y2232) );
  OA21x2_ASAP7_75t_R   g5038( .A1 (n407), .A2 (x2), .B (n3919), .Y (y2233) );
  NOR2x1_ASAP7_75t_R   g5039( .A (x5), .B (n1956), .Y (y2234) );
  OR3x1_ASAP7_75t_R    g5040( .A (x3), .B (x1), .C (x0), .Y (n5048) );
  INVx1_ASAP7_75t_R    g5041( .A (n5048), .Y (n5049) );
  AO21x1_ASAP7_75t_R   g5042( .A1 (n5049), .A2 (n15), .B (n131), .Y (y2235) );
  AO21x1_ASAP7_75t_R   g5043( .A1 (n218), .A2 (n22), .B (n3963), .Y (y2236) );
  AO21x1_ASAP7_75t_R   g5044( .A1 (y2079), .A2 (n3325), .B (n3386), .Y (y2237) );
  OR3x1_ASAP7_75t_R    g5045( .A (n1643), .B (n1644), .C (x0), .Y (y2239) );
  NAND2x1_ASAP7_75t_R  g5046( .A (y2079), .B (n3040), .Y (n5054) );
  INVx1_ASAP7_75t_R    g5047( .A (n5054), .Y (n5055) );
  OR3x1_ASAP7_75t_R    g5048( .A (n325), .B (y2079), .C (n12), .Y (n5056) );
  INVx1_ASAP7_75t_R    g5049( .A (n5056), .Y (n5057) );
  AO21x1_ASAP7_75t_R   g5050( .A1 (n348), .A2 (n5055), .B (n5057), .Y (y2240) );
  AO21x1_ASAP7_75t_R   g5051( .A1 (n1062), .A2 (n316), .B (x4), .Y (n5059) );
  NAND2x1_ASAP7_75t_R  g5052( .A (n5059), .B (n4520), .Y (y2241) );
  AO21x1_ASAP7_75t_R   g5053( .A1 (n17), .A2 (x4), .B (x0), .Y (n5061) );
  AND2x2_ASAP7_75t_R   g5054( .A (n556), .B (n5061), .Y (y2242) );
  AO32x1_ASAP7_75t_R   g5055( .A1 (n17), .A2 (n310), .A3 (n23), .B1 (x3), .B2 (y1281), .Y (y2243) );
  AND3x1_ASAP7_75t_R   g5056( .A (n72), .B (n137), .C (x5), .Y (n5064) );
  NAND2x1_ASAP7_75t_R  g5057( .A (x4), .B (n5064), .Y (n5065) );
  AO21x1_ASAP7_75t_R   g5058( .A1 (n3000), .A2 (n672), .B (n45), .Y (n5066) );
  AND2x2_ASAP7_75t_R   g5059( .A (n5065), .B (n5066), .Y (y2244) );
  NOR2x1_ASAP7_75t_R   g5060( .A (n481), .B (n375), .Y (y2245) );
  AO21x1_ASAP7_75t_R   g5061( .A1 (n301), .A2 (n299), .B (n989), .Y (y2246) );
  OA21x2_ASAP7_75t_R   g5062( .A1 (n1646), .A2 (n3035), .B (n2532), .Y (y2247) );
  AND2x2_ASAP7_75t_R   g5063( .A (n463), .B (n938), .Y (y2248) );
  INVx1_ASAP7_75t_R    g5064( .A (n3638), .Y (n5072) );
  OA21x2_ASAP7_75t_R   g5065( .A1 (n5072), .A2 (n4495), .B (n3286), .Y (y2249) );
  AO21x1_ASAP7_75t_R   g5066( .A1 (n1921), .A2 (y2079), .B (n977), .Y (y2251) );
  AND3x1_ASAP7_75t_R   g5067( .A (y855), .B (n228), .C (y2079), .Y (y2252) );
  AND2x2_ASAP7_75t_R   g5068( .A (n382), .B (n652), .Y (n5076) );
  NOR2x1_ASAP7_75t_R   g5069( .A (x5), .B (n5076), .Y (n5077) );
  AO21x1_ASAP7_75t_R   g5070( .A1 (n17), .A2 (n914), .B (n5077), .Y (y2253) );
  AO21x1_ASAP7_75t_R   g5071( .A1 (n52), .A2 (x0), .B (n716), .Y (y2254) );
  INVx1_ASAP7_75t_R    g5072( .A (n4723), .Y (n5080) );
  OR3x1_ASAP7_75t_R    g5073( .A (n363), .B (n22), .C (x3), .Y (n5081) );
  OA21x2_ASAP7_75t_R   g5074( .A1 (n5080), .A2 (n291), .B (n5081), .Y (y2255) );
  AND2x2_ASAP7_75t_R   g5075( .A (y1873), .B (n1265), .Y (y2256) );
  AO21x1_ASAP7_75t_R   g5076( .A1 (x4), .A2 (n17), .B (n97), .Y (n5084) );
  AO21x1_ASAP7_75t_R   g5077( .A1 (n15), .A2 (x5), .B (n22), .Y (n5085) );
  INVx1_ASAP7_75t_R    g5078( .A (n5085), .Y (n5086) );
  NAND2x1_ASAP7_75t_R  g5079( .A (n17), .B (n5086), .Y (n5087) );
  NAND2x1_ASAP7_75t_R  g5080( .A (n5084), .B (n5087), .Y (n5088) );
  OR3x1_ASAP7_75t_R    g5081( .A (n5088), .B (n3568), .C (n3443), .Y (y2257) );
  AO21x1_ASAP7_75t_R   g5082( .A1 (n22), .A2 (y2079), .B (x2), .Y (n5090) );
  NAND2x1_ASAP7_75t_R  g5083( .A (x3), .B (n5090), .Y (n5091) );
  AND2x2_ASAP7_75t_R   g5084( .A (n5091), .B (n4108), .Y (y2258) );
  OA21x2_ASAP7_75t_R   g5085( .A1 (n1851), .A2 (n671), .B (y2068), .Y (y2260) );
  INVx1_ASAP7_75t_R    g5086( .A (n3294), .Y (n5094) );
  AND3x1_ASAP7_75t_R   g5087( .A (n3943), .B (n5094), .C (n388), .Y (n5095) );
  INVx1_ASAP7_75t_R    g5088( .A (n5095), .Y (y2261) );
  OR3x1_ASAP7_75t_R    g5089( .A (n337), .B (y2079), .C (x2), .Y (n5097) );
  INVx1_ASAP7_75t_R    g5090( .A (n5097), .Y (n5098) );
  AND3x1_ASAP7_75t_R   g5091( .A (n406), .B (n632), .C (x2), .Y (n5099) );
  AO21x1_ASAP7_75t_R   g5092( .A1 (n5098), .A2 (n22), .B (n5099), .Y (y2262) );
  NOR2x1_ASAP7_75t_R   g5093( .A (x0), .B (n753), .Y (n5101) );
  AO21x1_ASAP7_75t_R   g5094( .A1 (n2508), .A2 (x1), .B (n5101), .Y (y2263) );
  OR3x1_ASAP7_75t_R    g5095( .A (n537), .B (x5), .C (x3), .Y (n5103) );
  AND2x2_ASAP7_75t_R   g5096( .A (y1777), .B (n5103), .Y (y2264) );
  INVx1_ASAP7_75t_R    g5097( .A (n2047), .Y (n5105) );
  OR3x1_ASAP7_75t_R    g5098( .A (n2169), .B (n363), .C (n128), .Y (n5106) );
  AND2x2_ASAP7_75t_R   g5099( .A (n5105), .B (n5106), .Y (y2265) );
  INVx1_ASAP7_75t_R    g5100( .A (n3207), .Y (n5108) );
  AO21x1_ASAP7_75t_R   g5101( .A1 (n740), .A2 (n17), .B (n3905), .Y (n5109) );
  OA21x2_ASAP7_75t_R   g5102( .A1 (n3298), .A2 (n5108), .B (n5109), .Y (y2266) );
  INVx1_ASAP7_75t_R    g5103( .A (n4635), .Y (n5111) );
  AO21x1_ASAP7_75t_R   g5104( .A1 (n5111), .A2 (y2079), .B (n3386), .Y (y2267) );
  AND3x1_ASAP7_75t_R   g5105( .A (n3109), .B (n2573), .C (n348), .Y (y2268) );
  AO21x1_ASAP7_75t_R   g5106( .A1 (n546), .A2 (n497), .B (n12), .Y (n5114) );
  OA21x2_ASAP7_75t_R   g5107( .A1 (x0), .A2 (n1992), .B (n5114), .Y (y2269) );
  AO21x1_ASAP7_75t_R   g5108( .A1 (x4), .A2 (x3), .B (n15), .Y (n5116) );
  INVx1_ASAP7_75t_R    g5109( .A (n5116), .Y (n5117) );
  OA21x2_ASAP7_75t_R   g5110( .A1 (n5117), .A2 (n3310), .B (y2079), .Y (y2270) );
  NOR2x1_ASAP7_75t_R   g5111( .A (n444), .B (n1927), .Y (y2271) );
  AND2x2_ASAP7_75t_R   g5112( .A (n4864), .B (n17), .Y (n5120) );
  AO21x1_ASAP7_75t_R   g5113( .A1 (y3758), .A2 (x3), .B (n5120), .Y (y2272) );
  AND2x2_ASAP7_75t_R   g5114( .A (n1480), .B (n747), .Y (y2273) );
  AO32x1_ASAP7_75t_R   g5115( .A1 (n700), .A2 (n3498), .A3 (n144), .B1 (n219), .B2 (n1215), .Y (y2275) );
  OR3x1_ASAP7_75t_R    g5116( .A (n403), .B (y2079), .C (n15), .Y (n5124) );
  INVx1_ASAP7_75t_R    g5117( .A (n5124), .Y (n5125) );
  AO21x1_ASAP7_75t_R   g5118( .A1 (n3565), .A2 (n3285), .B (n5125), .Y (y2276) );
  AO21x1_ASAP7_75t_R   g5119( .A1 (n17), .A2 (x2), .B (x4), .Y (n5127) );
  AO21x1_ASAP7_75t_R   g5120( .A1 (n15), .A2 (x3), .B (n22), .Y (n5128) );
  NAND2x1_ASAP7_75t_R  g5121( .A (n5127), .B (n5128), .Y (n5129) );
  AND2x2_ASAP7_75t_R   g5122( .A (n5129), .B (y3377), .Y (y2277) );
  AND2x2_ASAP7_75t_R   g5123( .A (n3625), .B (n4674), .Y (y2278) );
  AO21x1_ASAP7_75t_R   g5124( .A1 (n645), .A2 (n3327), .B (n22), .Y (n5132) );
  OA21x2_ASAP7_75t_R   g5125( .A1 (x4), .A2 (n323), .B (n5132), .Y (y2279) );
  AO21x1_ASAP7_75t_R   g5126( .A1 (n3192), .A2 (n22), .B (n363), .Y (y2281) );
  AND2x2_ASAP7_75t_R   g5127( .A (n3128), .B (y2079), .Y (y2282) );
  AO21x1_ASAP7_75t_R   g5128( .A1 (n64), .A2 (n2158), .B (n854), .Y (y2283) );
  OR3x1_ASAP7_75t_R    g5129( .A (n628), .B (n3263), .C (n3279), .Y (y2284) );
  AO21x1_ASAP7_75t_R   g5130( .A1 (n421), .A2 (n299), .B (n4523), .Y (y2285) );
  AND3x1_ASAP7_75t_R   g5131( .A (n1196), .B (y1894), .C (n471), .Y (y2286) );
  OR3x1_ASAP7_75t_R    g5132( .A (n518), .B (n16), .C (n12), .Y (n5140) );
  INVx1_ASAP7_75t_R    g5133( .A (n5140), .Y (n5141) );
  AO21x1_ASAP7_75t_R   g5134( .A1 (y2079), .A2 (n1007), .B (n5141), .Y (y2287) );
  AO21x1_ASAP7_75t_R   g5135( .A1 (n401), .A2 (n3565), .B (n756), .Y (n5143) );
  AND2x2_ASAP7_75t_R   g5136( .A (n4241), .B (n5143), .Y (y2288) );
  NAND2x1_ASAP7_75t_R  g5137( .A (n22), .B (n1092), .Y (n5145) );
  OA21x2_ASAP7_75t_R   g5138( .A1 (n590), .A2 (n22), .B (n5145), .Y (y2289) );
  INVx1_ASAP7_75t_R    g5139( .A (n4768), .Y (y2643) );
  OR3x1_ASAP7_75t_R    g5140( .A (n3027), .B (x5), .C (x3), .Y (n5148) );
  AND2x2_ASAP7_75t_R   g5141( .A (y2643), .B (n5148), .Y (y2290) );
  AO21x1_ASAP7_75t_R   g5142( .A1 (n527), .A2 (n765), .B (n1779), .Y (y2291) );
  AO21x1_ASAP7_75t_R   g5143( .A1 (n76), .A2 (x4), .B (x5), .Y (n5151) );
  INVx1_ASAP7_75t_R    g5144( .A (n5151), .Y (y2292) );
  AO21x1_ASAP7_75t_R   g5145( .A1 (n510), .A2 (n343), .B (x1), .Y (n5153) );
  AND2x2_ASAP7_75t_R   g5146( .A (n5153), .B (n1272), .Y (y2293) );
  AO21x1_ASAP7_75t_R   g5147( .A1 (y2079), .A2 (n507), .B (n914), .Y (y2483) );
  AND2x2_ASAP7_75t_R   g5148( .A (n1863), .B (y2483), .Y (y2294) );
  OA21x2_ASAP7_75t_R   g5149( .A1 (n73), .A2 (n121), .B (n118), .Y (y2295) );
  OR3x1_ASAP7_75t_R    g5150( .A (n5117), .B (y2079), .C (n3310), .Y (y2296) );
  INVx1_ASAP7_75t_R    g5151( .A (n4467), .Y (n5159) );
  AND2x2_ASAP7_75t_R   g5152( .A (n3804), .B (n5159), .Y (y2421) );
  INVx1_ASAP7_75t_R    g5153( .A (y2421), .Y (n5161) );
  AND3x1_ASAP7_75t_R   g5154( .A (n5161), .B (y1267), .C (n4070), .Y (y2297) );
  NAND2x1_ASAP7_75t_R  g5155( .A (x5), .B (n374), .Y (y2298) );
  AO21x1_ASAP7_75t_R   g5156( .A1 (x3), .A2 (n537), .B (n4920), .Y (n5164) );
  AO32x1_ASAP7_75t_R   g5157( .A1 (n1319), .A2 (n4289), .A3 (n58), .B1 (y2079), .B2 (n5164), .Y (y2299) );
  AO21x1_ASAP7_75t_R   g5158( .A1 (n28), .A2 (x3), .B (n2063), .Y (n5166) );
  INVx1_ASAP7_75t_R    g5159( .A (n5166), .Y (n5167) );
  AO21x1_ASAP7_75t_R   g5160( .A1 (x3), .A2 (n1775), .B (n5167), .Y (y2300) );
  AND2x2_ASAP7_75t_R   g5161( .A (y2737), .B (n1111), .Y (y2301) );
  NAND2x1_ASAP7_75t_R  g5162( .A (n295), .B (n125), .Y (y2716) );
  AND2x2_ASAP7_75t_R   g5163( .A (y2716), .B (n1370), .Y (y2302) );
  AO21x1_ASAP7_75t_R   g5164( .A1 (n474), .A2 (n17), .B (n628), .Y (y2303) );
  AND3x1_ASAP7_75t_R   g5165( .A (x3), .B (x2), .C (x4), .Y (n5173) );
  OR3x1_ASAP7_75t_R    g5166( .A (n3316), .B (n5173), .C (n81), .Y (n5174) );
  NOR2x1_ASAP7_75t_R   g5167( .A (x5), .B (n5174), .Y (y2304) );
  AO21x1_ASAP7_75t_R   g5168( .A1 (y2079), .A2 (x2), .B (n17), .Y (n5176) );
  INVx1_ASAP7_75t_R    g5169( .A (n5176), .Y (n5177) );
  NAND2x1_ASAP7_75t_R  g5170( .A (n22), .B (n5177), .Y (n5178) );
  INVx1_ASAP7_75t_R    g5171( .A (n4180), .Y (n5179) );
  AND3x1_ASAP7_75t_R   g5172( .A (n5178), .B (n5179), .C (n556), .Y (y2306) );
  INVx1_ASAP7_75t_R    g5173( .A (n3992), .Y (n5181) );
  OA21x2_ASAP7_75t_R   g5174( .A1 (n3132), .A2 (n22), .B (n5181), .Y (y2307) );
  OR3x1_ASAP7_75t_R    g5175( .A (n368), .B (x4), .C (x0), .Y (n5183) );
  AO21x1_ASAP7_75t_R   g5176( .A1 (n12), .A2 (y2079), .B (n4250), .Y (n5184) );
  AND2x2_ASAP7_75t_R   g5177( .A (n5183), .B (n5184), .Y (y2308) );
  AND3x1_ASAP7_75t_R   g5178( .A (n455), .B (n366), .C (x2), .Y (n5186) );
  AO21x1_ASAP7_75t_R   g5179( .A1 (n15), .A2 (n4099), .B (n5186), .Y (y2309) );
  OA21x2_ASAP7_75t_R   g5180( .A1 (n3298), .A2 (n5108), .B (n3943), .Y (y2310) );
  AO32x1_ASAP7_75t_R   g5181( .A1 (n17), .A2 (n3567), .A3 (x5), .B1 (n4916), .B2 (n556), .Y (y2311) );
  NOR2x1_ASAP7_75t_R   g5182( .A (x5), .B (n1911), .Y (n5190) );
  AO21x1_ASAP7_75t_R   g5183( .A1 (n5190), .A2 (y9), .B (n1778), .Y (y2312) );
  AO21x1_ASAP7_75t_R   g5184( .A1 (n3365), .A2 (n970), .B (n1948), .Y (y2313) );
  AND2x2_ASAP7_75t_R   g5185( .A (n1300), .B (y2079), .Y (n5193) );
  OR3x1_ASAP7_75t_R    g5186( .A (n5193), .B (n503), .C (n537), .Y (y2314) );
  AO21x1_ASAP7_75t_R   g5187( .A1 (n466), .A2 (y2079), .B (n58), .Y (y2315) );
  AO21x1_ASAP7_75t_R   g5188( .A1 (n1340), .A2 (n497), .B (x0), .Y (y2374) );
  NAND2x1_ASAP7_75t_R  g5189( .A (y2374), .B (n2092), .Y (y2316) );
  OA21x2_ASAP7_75t_R   g5190( .A1 (x0), .A2 (n1173), .B (n1046), .Y (y2317) );
  AND2x2_ASAP7_75t_R   g5191( .A (n3987), .B (y1359), .Y (y2318) );
  NAND2x1_ASAP7_75t_R  g5192( .A (n3024), .B (n3083), .Y (y2319) );
  AO21x1_ASAP7_75t_R   g5193( .A1 (n334), .A2 (x5), .B (n337), .Y (n5201) );
  INVx1_ASAP7_75t_R    g5194( .A (n5201), .Y (y2320) );
  AOI21x1_ASAP7_75t_R  g5195( .A1 (n763), .A2 (n1590), .B (n2927), .Y (y2321) );
  AND2x2_ASAP7_75t_R   g5196( .A (n4643), .B (y3132), .Y (y2322) );
  AND3x1_ASAP7_75t_R   g5197( .A (n299), .B (n1166), .C (y2079), .Y (y2323) );
  AO21x1_ASAP7_75t_R   g5198( .A1 (y2079), .A2 (n3121), .B (n4349), .Y (y2324) );
  AND2x2_ASAP7_75t_R   g5199( .A (n4129), .B (y3527), .Y (y2325) );
  AO21x1_ASAP7_75t_R   g5200( .A1 (n29), .A2 (n16), .B (n957), .Y (y2326) );
  AND2x2_ASAP7_75t_R   g5201( .A (n125), .B (n84), .Y (n5209) );
  INVx1_ASAP7_75t_R    g5202( .A (n5209), .Y (n5210) );
  NOR2x1_ASAP7_75t_R   g5203( .A (n1676), .B (n5210), .Y (y2327) );
  AO21x1_ASAP7_75t_R   g5204( .A1 (x3), .A2 (x5), .B (n15), .Y (n5212) );
  NAND2x1_ASAP7_75t_R  g5205( .A (x3), .B (n3819), .Y (n5213) );
  INVx1_ASAP7_75t_R    g5206( .A (n5213), .Y (n5214) );
  AO21x1_ASAP7_75t_R   g5207( .A1 (n660), .A2 (n5212), .B (n5214), .Y (n5215) );
  AND2x2_ASAP7_75t_R   g5208( .A (n5215), .B (n3000), .Y (y2328) );
  AO21x1_ASAP7_75t_R   g5209( .A1 (n388), .A2 (n16), .B (x0), .Y (n5217) );
  OA21x2_ASAP7_75t_R   g5210( .A1 (n1907), .A2 (n5217), .B (n919), .Y (y2329) );
  AND3x1_ASAP7_75t_R   g5211( .A (n757), .B (n72), .C (n290), .Y (y2330) );
  NOR2x1_ASAP7_75t_R   g5212( .A (x5), .B (n4649), .Y (y2331) );
  AO32x1_ASAP7_75t_R   g5213( .A1 (n312), .A2 (n1426), .A3 (n1469), .B1 (x0), .B2 (n1643), .Y (y2332) );
  NOR2x1_ASAP7_75t_R   g5214( .A (n3376), .B (n139), .Y (y2333) );
  AND2x2_ASAP7_75t_R   g5215( .A (n463), .B (n1077), .Y (y2334) );
  AO21x1_ASAP7_75t_R   g5216( .A1 (x5), .A2 (x4), .B (n76), .Y (n5224) );
  INVx1_ASAP7_75t_R    g5217( .A (n5224), .Y (y2335) );
  AND3x1_ASAP7_75t_R   g5218( .A (n3387), .B (n3128), .C (y2079), .Y (y2336) );
  AO21x1_ASAP7_75t_R   g5219( .A1 (n17), .A2 (n22), .B (n15), .Y (n5227) );
  NAND2x1_ASAP7_75t_R  g5220( .A (n3526), .B (n5227), .Y (n5228) );
  AND2x2_ASAP7_75t_R   g5221( .A (n5228), .B (y2079), .Y (n5229) );
  AO21x1_ASAP7_75t_R   g5222( .A1 (n3493), .A2 (n29), .B (n5229), .Y (y2337) );
  AO21x1_ASAP7_75t_R   g5223( .A1 (n4375), .A2 (y2079), .B (n337), .Y (y2338) );
  AO21x1_ASAP7_75t_R   g5224( .A1 (n1215), .A2 (x0), .B (n2001), .Y (y2339) );
  INVx1_ASAP7_75t_R    g5225( .A (n591), .Y (n5233) );
  AO21x1_ASAP7_75t_R   g5226( .A1 (y435), .A2 (n5233), .B (n1959), .Y (y2340) );
  INVx1_ASAP7_75t_R    g5227( .A (n3315), .Y (n5235) );
  OR3x1_ASAP7_75t_R    g5228( .A (x4), .B (x3), .C (x2), .Y (n5236) );
  INVx1_ASAP7_75t_R    g5229( .A (n5236), .Y (n5237) );
  AO21x1_ASAP7_75t_R   g5230( .A1 (y2079), .A2 (n5235), .B (n5237), .Y (y2341) );
  AO21x1_ASAP7_75t_R   g5231( .A1 (n77), .A2 (x5), .B (n3447), .Y (n5239) );
  AO21x1_ASAP7_75t_R   g5232( .A1 (n5239), .A2 (n1572), .B (n529), .Y (y2342) );
  AND2x2_ASAP7_75t_R   g5233( .A (n1046), .B (n1272), .Y (y2343) );
  AND3x1_ASAP7_75t_R   g5234( .A (n189), .B (n572), .C (n369), .Y (y2344) );
  AO21x1_ASAP7_75t_R   g5235( .A1 (n22), .A2 (n17), .B (x2), .Y (n5243) );
  AND2x2_ASAP7_75t_R   g5236( .A (n382), .B (n5243), .Y (n5244) );
  NOR2x1_ASAP7_75t_R   g5237( .A (x5), .B (n5244), .Y (n5245) );
  AO21x1_ASAP7_75t_R   g5238( .A1 (n22), .A2 (n421), .B (n5245), .Y (y2345) );
  AND3x1_ASAP7_75t_R   g5239( .A (n28), .B (n84), .C (n125), .Y (n5247) );
  OR3x1_ASAP7_75t_R    g5240( .A (n399), .B (n389), .C (n5247), .Y (y2346) );
  INVx1_ASAP7_75t_R    g5241( .A (n3109), .Y (y2347) );
  NAND2x1_ASAP7_75t_R  g5242( .A (n388), .B (n360), .Y (n5250) );
  AND3x1_ASAP7_75t_R   g5243( .A (n369), .B (n388), .C (n15), .Y (n5251) );
  AO21x1_ASAP7_75t_R   g5244( .A1 (n5250), .A2 (x2), .B (n5251), .Y (y2348) );
  AO21x1_ASAP7_75t_R   g5245( .A1 (n700), .A2 (n22), .B (n363), .Y (n5253) );
  AO21x1_ASAP7_75t_R   g5246( .A1 (n533), .A2 (n5253), .B (n537), .Y (y2349) );
  AND2x2_ASAP7_75t_R   g5247( .A (n1851), .B (n463), .Y (y2350) );
  AO21x1_ASAP7_75t_R   g5248( .A1 (n22), .A2 (x2), .B (x5), .Y (n5256) );
  NOR2x1_ASAP7_75t_R   g5249( .A (n17), .B (n5256), .Y (n5257) );
  AO21x1_ASAP7_75t_R   g5250( .A1 (n17), .A2 (n3124), .B (n5257), .Y (y2351) );
  OR3x1_ASAP7_75t_R    g5251( .A (y3758), .B (n12), .C (n437), .Y (n5259) );
  OAI21x1_ASAP7_75t_R  g5252( .A1 (n396), .A2 (n580), .B (n5259), .Y (y2352) );
  AO21x1_ASAP7_75t_R   g5253( .A1 (n2116), .A2 (n244), .B (x5), .Y (n5261) );
  AND2x2_ASAP7_75t_R   g5254( .A (n5261), .B (n1405), .Y (y2353) );
  AND3x1_ASAP7_75t_R   g5255( .A (n465), .B (n466), .C (x0), .Y (y2354) );
  AND3x1_ASAP7_75t_R   g5256( .A (n3209), .B (n3469), .C (n632), .Y (y2355) );
  AO21x1_ASAP7_75t_R   g5257( .A1 (x1), .A2 (n2746), .B (n4784), .Y (y2356) );
  AO32x1_ASAP7_75t_R   g5258( .A1 (n144), .A2 (x2), .A3 (n700), .B1 (y1356), .B2 (n2463), .Y (n5266) );
  INVx1_ASAP7_75t_R    g5259( .A (n5266), .Y (y2357) );
  AO21x1_ASAP7_75t_R   g5260( .A1 (x5), .A2 (n3414), .B (n628), .Y (y2358) );
  AO21x1_ASAP7_75t_R   g5261( .A1 (n1927), .A2 (n17), .B (n4527), .Y (n5269) );
  AO21x1_ASAP7_75t_R   g5262( .A1 (x5), .A2 (n12), .B (n360), .Y (n5270) );
  INVx1_ASAP7_75t_R    g5263( .A (n5270), .Y (n5271) );
  AO21x1_ASAP7_75t_R   g5264( .A1 (n5269), .A2 (x0), .B (n5271), .Y (y2359) );
  AO21x1_ASAP7_75t_R   g5265( .A1 (n12), .A2 (n16), .B (n2576), .Y (n5273) );
  INVx1_ASAP7_75t_R    g5266( .A (n5273), .Y (n5274) );
  AO32x1_ASAP7_75t_R   g5267( .A1 (x2), .A2 (n3800), .A3 (n5274), .B1 (n15), .B2 (n5273), .Y (y2360) );
  OA21x2_ASAP7_75t_R   g5268( .A1 (n378), .A2 (n1265), .B (y3527), .Y (y2361) );
  AND2x2_ASAP7_75t_R   g5269( .A (n762), .B (n2885), .Y (y2362) );
  NAND2x1_ASAP7_75t_R  g5270( .A (n137), .B (n746), .Y (n5278) );
  AO21x1_ASAP7_75t_R   g5271( .A1 (n243), .A2 (n244), .B (n5278), .Y (n5279) );
  AND2x2_ASAP7_75t_R   g5272( .A (n4263), .B (n5279), .Y (y2363) );
  AO21x1_ASAP7_75t_R   g5273( .A1 (n3013), .A2 (n4619), .B (n418), .Y (n5281) );
  AND2x2_ASAP7_75t_R   g5274( .A (n5281), .B (n72), .Y (y2364) );
  AO21x1_ASAP7_75t_R   g5275( .A1 (n998), .A2 (n3203), .B (n2036), .Y (y2365) );
  OR3x1_ASAP7_75t_R    g5276( .A (n529), .B (n1158), .C (n2718), .Y (y2366) );
  AO21x1_ASAP7_75t_R   g5277( .A1 (n15), .A2 (x1), .B (y2079), .Y (n5285) );
  AO21x1_ASAP7_75t_R   g5278( .A1 (n64), .A2 (x0), .B (n5285), .Y (n5286) );
  OA21x2_ASAP7_75t_R   g5279( .A1 (n1596), .A2 (n4192), .B (n5286), .Y (y2367) );
  AND2x2_ASAP7_75t_R   g5280( .A (n2886), .B (x0), .Y (n5288) );
  AO21x1_ASAP7_75t_R   g5281( .A1 (x1), .A2 (n2210), .B (n5288), .Y (y2368) );
  AND2x2_ASAP7_75t_R   g5282( .A (y1267), .B (n4070), .Y (y2369) );
  OA21x2_ASAP7_75t_R   g5283( .A1 (n218), .A2 (y2079), .B (n2998), .Y (y2370) );
  OA21x2_ASAP7_75t_R   g5284( .A1 (n590), .A2 (n750), .B (n2182), .Y (y2371) );
  AO21x1_ASAP7_75t_R   g5285( .A1 (n1434), .A2 (n125), .B (x4), .Y (n5293) );
  OR3x1_ASAP7_75t_R    g5286( .A (n2718), .B (n388), .C (n425), .Y (n5294) );
  NAND2x1_ASAP7_75t_R  g5287( .A (n5293), .B (n5294), .Y (y2372) );
  AO21x1_ASAP7_75t_R   g5288( .A1 (y2079), .A2 (n22), .B (n15), .Y (n5296) );
  NAND2x1_ASAP7_75t_R  g5289( .A (x3), .B (n5296), .Y (n5297) );
  AND3x1_ASAP7_75t_R   g5290( .A (n5297), .B (n3013), .C (n3011), .Y (y2373) );
  AO21x1_ASAP7_75t_R   g5291( .A1 (n64), .A2 (n2158), .B (y2079), .Y (y2375) );
  OR3x1_ASAP7_75t_R    g5292( .A (n529), .B (n437), .C (n58), .Y (y2377) );
  AND2x2_ASAP7_75t_R   g5293( .A (n382), .B (y3377), .Y (y2378) );
  INVx1_ASAP7_75t_R    g5294( .A (n4469), .Y (y3676) );
  OR3x1_ASAP7_75t_R    g5295( .A (y2466), .B (n15), .C (n17), .Y (n5303) );
  INVx1_ASAP7_75t_R    g5296( .A (n5303), .Y (n5304) );
  OR3x1_ASAP7_75t_R    g5297( .A (y3676), .B (n5304), .C (n81), .Y (n5305) );
  NOR2x1_ASAP7_75t_R   g5298( .A (n518), .B (n5305), .Y (y2379) );
  AO21x1_ASAP7_75t_R   g5299( .A1 (n22), .A2 (n228), .B (n950), .Y (n5307) );
  OA21x2_ASAP7_75t_R   g5300( .A1 (n5307), .A2 (y863), .B (y2079), .Y (y2380) );
  AND2x2_ASAP7_75t_R   g5301( .A (y3397), .B (n455), .Y (y2381) );
  NAND2x1_ASAP7_75t_R  g5302( .A (n22), .B (n781), .Y (n5310) );
  OA21x2_ASAP7_75t_R   g5303( .A1 (n589), .A2 (n5310), .B (n2204), .Y (y2382) );
  AO21x1_ASAP7_75t_R   g5304( .A1 (n144), .A2 (n1646), .B (n2193), .Y (y2383) );
  AND2x2_ASAP7_75t_R   g5305( .A (n1176), .B (n463), .Y (y2384) );
  INVx1_ASAP7_75t_R    g5306( .A (n4495), .Y (n5314) );
  AND2x2_ASAP7_75t_R   g5307( .A (n3302), .B (n3377), .Y (y3366) );
  OA21x2_ASAP7_75t_R   g5308( .A1 (x5), .A2 (n5314), .B (y3366), .Y (y2385) );
  OA21x2_ASAP7_75t_R   g5309( .A1 (n421), .A2 (n4844), .B (n3944), .Y (y2386) );
  OR3x1_ASAP7_75t_R    g5310( .A (n128), .B (n12), .C (x5), .Y (n5318) );
  INVx1_ASAP7_75t_R    g5311( .A (n5318), .Y (y2387) );
  OR3x1_ASAP7_75t_R    g5312( .A (n51), .B (n12), .C (x3), .Y (n5320) );
  AO21x1_ASAP7_75t_R   g5313( .A1 (n2754), .A2 (n5320), .B (n13), .Y (y2388) );
  AO32x1_ASAP7_75t_R   g5314( .A1 (n360), .A2 (n290), .A3 (n5055), .B1 (n378), .B2 (n5054), .Y (y2390) );
  INVx1_ASAP7_75t_R    g5315( .A (n3918), .Y (n5323) );
  AND2x2_ASAP7_75t_R   g5316( .A (n3524), .B (n5323), .Y (n5324) );
  NOR2x1_ASAP7_75t_R   g5317( .A (n4768), .B (n5324), .Y (y2391) );
  OR3x1_ASAP7_75t_R    g5318( .A (n1248), .B (n58), .C (n128), .Y (n5326) );
  AND2x2_ASAP7_75t_R   g5319( .A (n5326), .B (n737), .Y (y2392) );
  AND3x1_ASAP7_75t_R   g5320( .A (n4142), .B (n77), .C (n556), .Y (y2394) );
  AO21x1_ASAP7_75t_R   g5321( .A1 (y2079), .A2 (x0), .B (n315), .Y (n5329) );
  OA21x2_ASAP7_75t_R   g5322( .A1 (n437), .A2 (n5329), .B (n2940), .Y (y2395) );
  AND3x1_ASAP7_75t_R   g5323( .A (n3250), .B (n22), .C (n17), .Y (n5331) );
  AO21x1_ASAP7_75t_R   g5324( .A1 (n401), .A2 (n3249), .B (n5331), .Y (y2396) );
  AO21x1_ASAP7_75t_R   g5325( .A1 (x4), .A2 (y2079), .B (n77), .Y (n5333) );
  AND2x2_ASAP7_75t_R   g5326( .A (n3549), .B (n5333), .Y (y2397) );
  AND2x2_ASAP7_75t_R   g5327( .A (n3374), .B (y2079), .Y (n5335) );
  AO21x1_ASAP7_75t_R   g5328( .A1 (n17), .A2 (n3124), .B (n5335), .Y (y2398) );
  AO21x1_ASAP7_75t_R   g5329( .A1 (n914), .A2 (n17), .B (y2079), .Y (n5337) );
  AND2x2_ASAP7_75t_R   g5330( .A (n4681), .B (n5337), .Y (y2399) );
  OR3x1_ASAP7_75t_R    g5331( .A (n3055), .B (n2994), .C (n628), .Y (y2400) );
  AND2x2_ASAP7_75t_R   g5332( .A (y109), .B (n546), .Y (y2401) );
  OA21x2_ASAP7_75t_R   g5333( .A1 (n2445), .A2 (n3365), .B (n2940), .Y (y2402) );
  AO21x1_ASAP7_75t_R   g5334( .A1 (n316), .A2 (n319), .B (n310), .Y (n5342) );
  OA21x2_ASAP7_75t_R   g5335( .A1 (n4360), .A2 (n4361), .B (n5342), .Y (y2403) );
  AO21x1_ASAP7_75t_R   g5336( .A1 (n3880), .A2 (n1125), .B (n529), .Y (y2404) );
  AND2x2_ASAP7_75t_R   g5337( .A (n401), .B (n299), .Y (n5345) );
  AO21x1_ASAP7_75t_R   g5338( .A1 (n5345), .A2 (y2079), .B (n4349), .Y (y2405) );
  OR3x1_ASAP7_75t_R    g5339( .A (n1158), .B (y2079), .C (n2994), .Y (y3427) );
  AND2x2_ASAP7_75t_R   g5340( .A (y3427), .B (n4508), .Y (y2406) );
  AO21x1_ASAP7_75t_R   g5341( .A1 (n285), .A2 (n287), .B (x2), .Y (n5349) );
  AND2x2_ASAP7_75t_R   g5342( .A (n4571), .B (n5349), .Y (y2407) );
  AND3x1_ASAP7_75t_R   g5343( .A (n128), .B (n12), .C (x3), .Y (n5351) );
  AO21x1_ASAP7_75t_R   g5344( .A1 (n129), .A2 (x0), .B (n5351), .Y (y2408) );
  AND2x2_ASAP7_75t_R   g5345( .A (n4945), .B (n2701), .Y (y2409) );
  NOR2x1_ASAP7_75t_R   g5346( .A (n17), .B (n537), .Y (n5354) );
  NAND2x1_ASAP7_75t_R  g5347( .A (n22), .B (n3646), .Y (n5355) );
  OA211x2_ASAP7_75t_R  g5348( .A1 (n1164), .A2 (n5354), .B (n5355), .C (y3852), .Y (y2410) );
  AO21x1_ASAP7_75t_R   g5349( .A1 (n671), .A2 (n15), .B (n76), .Y (n5357) );
  OA211x2_ASAP7_75t_R  g5350( .A1 (n22), .A2 (n5357), .B (n3655), .C (n2971), .Y (y2411) );
  AO21x1_ASAP7_75t_R   g5351( .A1 (y9), .A2 (n529), .B (n1083), .Y (y2412) );
  AO21x1_ASAP7_75t_R   g5352( .A1 (n529), .A2 (n1062), .B (n3025), .Y (y2413) );
  INVx1_ASAP7_75t_R    g5353( .A (n5008), .Y (y2414) );
  AO21x1_ASAP7_75t_R   g5354( .A1 (n22), .A2 (x3), .B (x5), .Y (n5362) );
  INVx1_ASAP7_75t_R    g5355( .A (n5362), .Y (n5363) );
  OA21x2_ASAP7_75t_R   g5356( .A1 (n218), .A2 (n5363), .B (n4647), .Y (y2415) );
  AO21x1_ASAP7_75t_R   g5357( .A1 (x2), .A2 (n978), .B (y772), .Y (y2416) );
  AO21x1_ASAP7_75t_R   g5358( .A1 (n455), .A2 (n757), .B (n1158), .Y (n5366) );
  AND2x2_ASAP7_75t_R   g5359( .A (n5366), .B (n72), .Y (y2417) );
  AO21x1_ASAP7_75t_R   g5360( .A1 (n1851), .A2 (n17), .B (n2843), .Y (n5368) );
  AND3x1_ASAP7_75t_R   g5361( .A (n5368), .B (n4559), .C (n556), .Y (y2418) );
  AND3x1_ASAP7_75t_R   g5362( .A (y3293), .B (n137), .C (n72), .Y (n5370) );
  AND2x2_ASAP7_75t_R   g5363( .A (n5370), .B (n3014), .Y (y2419) );
  AO21x1_ASAP7_75t_R   g5364( .A1 (n12), .A2 (n22), .B (n17), .Y (n5372) );
  INVx1_ASAP7_75t_R    g5365( .A (n5372), .Y (n5373) );
  OA33x2_ASAP7_75t_R   g5366( .A1 (n17), .A2 (n22), .A3 (y2079), .B1 (n368), .B2 (n5373), .B3 (n537), .Y (y2420) );
  AO21x1_ASAP7_75t_R   g5367( .A1 (y2196), .A2 (n348), .B (n4514), .Y (y2422) );
  AND3x1_ASAP7_75t_R   g5368( .A (y1903), .B (n4336), .C (n672), .Y (y2423) );
  AO21x1_ASAP7_75t_R   g5369( .A1 (n382), .A2 (x0), .B (n349), .Y (y2424) );
  AO21x1_ASAP7_75t_R   g5370( .A1 (n17), .A2 (n22), .B (n3636), .Y (n5378) );
  AOI21x1_ASAP7_75t_R  g5371( .A1 (n4495), .A2 (n5378), .B (n518), .Y (y2425) );
  OR3x1_ASAP7_75t_R    g5372( .A (n103), .B (n17), .C (x0), .Y (n5380) );
  INVx1_ASAP7_75t_R    g5373( .A (n5380), .Y (n5381) );
  NOR2x1_ASAP7_75t_R   g5374( .A (n12), .B (n105), .Y (n5382) );
  OR3x1_ASAP7_75t_R    g5375( .A (n5381), .B (n5382), .C (n128), .Y (y2426) );
  AND3x1_ASAP7_75t_R   g5376( .A (n1391), .B (n2407), .C (y2079), .Y (y2427) );
  INVx1_ASAP7_75t_R    g5377( .A (n5256), .Y (n5385) );
  AO21x1_ASAP7_75t_R   g5378( .A1 (n5385), .A2 (x3), .B (n337), .Y (y2428) );
  AND2x2_ASAP7_75t_R   g5379( .A (n380), .B (y1865), .Y (y2429) );
  OR3x1_ASAP7_75t_R    g5380( .A (n2147), .B (n791), .C (y2196), .Y (y2430) );
  AND2x2_ASAP7_75t_R   g5381( .A (y2727), .B (n632), .Y (y2431) );
  AO21x1_ASAP7_75t_R   g5382( .A1 (n15), .A2 (x4), .B (n211), .Y (n5390) );
  AO21x1_ASAP7_75t_R   g5383( .A1 (n5390), .A2 (y2079), .B (n337), .Y (y2433) );
  AO21x1_ASAP7_75t_R   g5384( .A1 (y9), .A2 (n29), .B (n1078), .Y (y2434) );
  AO21x1_ASAP7_75t_R   g5385( .A1 (x1), .A2 (x0), .B (n17), .Y (n5393) );
  OA21x2_ASAP7_75t_R   g5386( .A1 (n3937), .A2 (n1669), .B (n5393), .Y (y2435) );
  AO21x1_ASAP7_75t_R   g5387( .A1 (y2079), .A2 (n3128), .B (n3386), .Y (y2436) );
  AO21x1_ASAP7_75t_R   g5388( .A1 (n948), .A2 (y2079), .B (y863), .Y (y2904) );
  AND2x2_ASAP7_75t_R   g5389( .A (y2904), .B (n947), .Y (y2437) );
  AND3x1_ASAP7_75t_R   g5390( .A (n137), .B (n22), .C (y2079), .Y (n5398) );
  INVx1_ASAP7_75t_R    g5391( .A (n5398), .Y (n5399) );
  AND2x2_ASAP7_75t_R   g5392( .A (n5399), .B (y1388), .Y (y2438) );
  AO21x1_ASAP7_75t_R   g5393( .A1 (x0), .A2 (x4), .B (n17), .Y (n5401) );
  AND3x1_ASAP7_75t_R   g5394( .A (n290), .B (y1281), .C (n5401), .Y (y2439) );
  AND2x2_ASAP7_75t_R   g5395( .A (n3284), .B (x0), .Y (n5403) );
  OA21x2_ASAP7_75t_R   g5396( .A1 (n3112), .A2 (n5403), .B (n3256), .Y (y2440) );
  AO21x1_ASAP7_75t_R   g5397( .A1 (n129), .A2 (x0), .B (n2047), .Y (y2441) );
  INVx1_ASAP7_75t_R    g5398( .A (n647), .Y (y2443) );
  OA21x2_ASAP7_75t_R   g5399( .A1 (n4584), .A2 (n604), .B (n642), .Y (y2444) );
  OA21x2_ASAP7_75t_R   g5400( .A1 (n1215), .A2 (n315), .B (n219), .Y (y2445) );
  AO21x1_ASAP7_75t_R   g5401( .A1 (y2079), .A2 (x4), .B (n1150), .Y (y2446) );
  AO21x1_ASAP7_75t_R   g5402( .A1 (n125), .A2 (x4), .B (n3386), .Y (n5410) );
  INVx1_ASAP7_75t_R    g5403( .A (n5410), .Y (n5411) );
  AO21x1_ASAP7_75t_R   g5404( .A1 (n5411), .A2 (n3160), .B (n3129), .Y (y2447) );
  AO21x1_ASAP7_75t_R   g5405( .A1 (y2079), .A2 (n3143), .B (n337), .Y (n5413) );
  AND2x2_ASAP7_75t_R   g5406( .A (n5413), .B (n4374), .Y (y2448) );
  AND3x1_ASAP7_75t_R   g5407( .A (n4821), .B (n724), .C (y3377), .Y (y2449) );
  NAND2x1_ASAP7_75t_R  g5408( .A (n690), .B (n310), .Y (y2450) );
  AO21x1_ASAP7_75t_R   g5409( .A1 (n583), .A2 (n16), .B (n1529), .Y (n5417) );
  OA21x2_ASAP7_75t_R   g5410( .A1 (n15), .A2 (y873), .B (n5417), .Y (y2451) );
  AO21x1_ASAP7_75t_R   g5411( .A1 (n368), .A2 (n22), .B (x2), .Y (n5419) );
  OA21x2_ASAP7_75t_R   g5412( .A1 (y2068), .A2 (n15), .B (n5419), .Y (y2452) );
  NAND2x1_ASAP7_75t_R  g5413( .A (n1707), .B (n388), .Y (y2453) );
  AO21x1_ASAP7_75t_R   g5414( .A1 (n299), .A2 (n310), .B (x1), .Y (n5422) );
  INVx1_ASAP7_75t_R    g5415( .A (n5422), .Y (n5423) );
  AO21x1_ASAP7_75t_R   g5416( .A1 (x4), .A2 (n12), .B (n776), .Y (n5424) );
  INVx1_ASAP7_75t_R    g5417( .A (n5424), .Y (n5425) );
  OR3x1_ASAP7_75t_R    g5418( .A (n5423), .B (n5425), .C (n529), .Y (y2454) );
  INVx1_ASAP7_75t_R    g5419( .A (n4109), .Y (n5427) );
  OR3x1_ASAP7_75t_R    g5420( .A (n5427), .B (n3263), .C (n1269), .Y (y2455) );
  INVx1_ASAP7_75t_R    g5421( .A (n906), .Y (y2456) );
  NOR2x1_ASAP7_75t_R   g5422( .A (x5), .B (n4465), .Y (y2457) );
  AND3x1_ASAP7_75t_R   g5423( .A (y3293), .B (n457), .C (x0), .Y (y2458) );
  AND2x2_ASAP7_75t_R   g5424( .A (y1693), .B (n3884), .Y (y2459) );
  AND3x1_ASAP7_75t_R   g5425( .A (n28), .B (n299), .C (n16), .Y (n5433) );
  NOR2x1_ASAP7_75t_R   g5426( .A (n481), .B (n5433), .Y (y2460) );
  AO21x1_ASAP7_75t_R   g5427( .A1 (n299), .A2 (y2079), .B (n17), .Y (n5435) );
  OA21x2_ASAP7_75t_R   g5428( .A1 (x3), .A2 (n474), .B (n5435), .Y (y2461) );
  AO21x1_ASAP7_75t_R   g5429( .A1 (n3738), .A2 (y6), .B (n2107), .Y (y2462) );
  INVx1_ASAP7_75t_R    g5430( .A (n3944), .Y (n5438) );
  NOR2x1_ASAP7_75t_R   g5431( .A (n5438), .B (n4910), .Y (y2463) );
  AO21x1_ASAP7_75t_R   g5432( .A1 (n17), .A2 (x2), .B (n518), .Y (n5440) );
  INVx1_ASAP7_75t_R    g5433( .A (n5440), .Y (n5441) );
  OR3x1_ASAP7_75t_R    g5434( .A (n856), .B (n22), .C (x3), .Y (n5442) );
  INVx1_ASAP7_75t_R    g5435( .A (n5442), .Y (n5443) );
  AO21x1_ASAP7_75t_R   g5436( .A1 (n290), .A2 (n5441), .B (n5443), .Y (y2465) );
  AO21x1_ASAP7_75t_R   g5437( .A1 (n2776), .A2 (n3354), .B (n4448), .Y (y2467) );
  AND2x2_ASAP7_75t_R   g5438( .A (n2998), .B (x5), .Y (n5446) );
  OA21x2_ASAP7_75t_R   g5439( .A1 (n217), .A2 (n5446), .B (n3002), .Y (y2468) );
  AO21x1_ASAP7_75t_R   g5440( .A1 (y104), .A2 (n1997), .B (n139), .Y (y2469) );
  AO21x1_ASAP7_75t_R   g5441( .A1 (x3), .A2 (n22), .B (n2971), .Y (n5449) );
  AND2x2_ASAP7_75t_R   g5442( .A (n5449), .B (n4695), .Y (y2470) );
  INVx1_ASAP7_75t_R    g5443( .A (n4317), .Y (n5451) );
  OA21x2_ASAP7_75t_R   g5444( .A1 (n5451), .A2 (y2740), .B (n1265), .Y (y2471) );
  AO21x1_ASAP7_75t_R   g5445( .A1 (y2079), .A2 (n4371), .B (n4529), .Y (y2472) );
  OA22x2_ASAP7_75t_R   g5446( .A1 (n756), .A2 (n3776), .B1 (n3294), .B2 (n4903), .Y (y2473) );
  AO32x1_ASAP7_75t_R   g5447( .A1 (n348), .A2 (y3852), .A3 (n3109), .B1 (n481), .B2 (n382), .Y (y2474) );
  OR3x1_ASAP7_75t_R    g5448( .A (n1004), .B (n478), .C (n143), .Y (y2475) );
  NOR2x1_ASAP7_75t_R   g5449( .A (n3608), .B (n4486), .Y (n5457) );
  OA21x2_ASAP7_75t_R   g5450( .A1 (n15), .A2 (y2443), .B (n5457), .Y (y2476) );
  OA33x2_ASAP7_75t_R   g5451( .A1 (n15), .A2 (x4), .A3 (n421), .B1 (n1269), .B2 (n3568), .B3 (n1158), .Y (y2477) );
  AND3x1_ASAP7_75t_R   g5452( .A (n3261), .B (n3327), .C (n645), .Y (y2478) );
  AND2x2_ASAP7_75t_R   g5453( .A (n1319), .B (y2079), .Y (n5461) );
  AO21x1_ASAP7_75t_R   g5454( .A1 (n5461), .A2 (n189), .B (n638), .Y (y2479) );
  OR3x1_ASAP7_75t_R    g5455( .A (n17), .B (y2079), .C (x0), .Y (n5463) );
  AO21x1_ASAP7_75t_R   g5456( .A1 (n3256), .A2 (n5463), .B (n306), .Y (y2480) );
  AO21x1_ASAP7_75t_R   g5457( .A1 (n72), .A2 (n137), .B (x4), .Y (n5465) );
  INVx1_ASAP7_75t_R    g5458( .A (n5465), .Y (n5466) );
  AO21x1_ASAP7_75t_R   g5459( .A1 (n72), .A2 (n529), .B (n5466), .Y (y2481) );
  AOI22x1_ASAP7_75t_R  g5460( .A1 (n3857), .A2 (x5), .B1 (n3776), .B2 (n15), .Y (y2484) );
  AO21x1_ASAP7_75t_R   g5461( .A1 (x5), .A2 (n914), .B (y2172), .Y (y2485) );
  OA21x2_ASAP7_75t_R   g5462( .A1 (x0), .A2 (n464), .B (n3380), .Y (y2486) );
  INVx1_ASAP7_75t_R    g5463( .A (n4057), .Y (n5471) );
  AO32x1_ASAP7_75t_R   g5464( .A1 (n17), .A2 (n5085), .A3 (n5471), .B1 (x3), .B2 (n4057), .Y (y2487) );
  AO21x1_ASAP7_75t_R   g5465( .A1 (n29), .A2 (n77), .B (n4575), .Y (y2488) );
  OA21x2_ASAP7_75t_R   g5466( .A1 (y772), .A2 (n1636), .B (n2701), .Y (y2489) );
  OA21x2_ASAP7_75t_R   g5467( .A1 (n2455), .A2 (n2315), .B (n2524), .Y (y2491) );
  AND3x1_ASAP7_75t_R   g5468( .A (n137), .B (y2079), .C (n22), .Y (n5476) );
  INVx1_ASAP7_75t_R    g5469( .A (y3397), .Y (n5477) );
  NOR2x1_ASAP7_75t_R   g5470( .A (n5476), .B (n5477), .Y (y2492) );
  OR3x1_ASAP7_75t_R    g5471( .A (n1032), .B (n3519), .C (x4), .Y (n5479) );
  AND2x2_ASAP7_75t_R   g5472( .A (n5479), .B (y1903), .Y (y2493) );
  OA21x2_ASAP7_75t_R   g5473( .A1 (n914), .A2 (n403), .B (n369), .Y (y2494) );
  AND3x1_ASAP7_75t_R   g5474( .A (n757), .B (n290), .C (n4495), .Y (n5482) );
  INVx1_ASAP7_75t_R    g5475( .A (n5482), .Y (n5483) );
  AO21x1_ASAP7_75t_R   g5476( .A1 (n290), .A2 (y2079), .B (n4495), .Y (n5484) );
  AND2x2_ASAP7_75t_R   g5477( .A (n5483), .B (n5484), .Y (y2495) );
  OA21x2_ASAP7_75t_R   g5478( .A1 (n3963), .A2 (n22), .B (n3655), .Y (y2496) );
  OA22x2_ASAP7_75t_R   g5479( .A1 (n4526), .A2 (n5314), .B1 (n5466), .B2 (n3960), .Y (y2497) );
  OR3x1_ASAP7_75t_R    g5480( .A (n4584), .B (n1817), .C (n145), .Y (y2499) );
  OR3x1_ASAP7_75t_R    g5481( .A (y1081), .B (n182), .C (n787), .Y (y2501) );
  NOR2x1_ASAP7_75t_R   g5482( .A (n518), .B (n1182), .Y (y2502) );
  OA21x2_ASAP7_75t_R   g5483( .A1 (n4116), .A2 (n3502), .B (n3648), .Y (y2503) );
  AO21x1_ASAP7_75t_R   g5484( .A1 (x5), .A2 (n5076), .B (n5077), .Y (y3598) );
  INVx1_ASAP7_75t_R    g5485( .A (n3189), .Y (n5493) );
  AND2x2_ASAP7_75t_R   g5486( .A (y3598), .B (n5493), .Y (y2504) );
  NAND2x1_ASAP7_75t_R  g5487( .A (n1092), .B (n3404), .Y (n5495) );
  AND2x2_ASAP7_75t_R   g5488( .A (n5495), .B (y1281), .Y (y2505) );
  INVx1_ASAP7_75t_R    g5489( .A (n4200), .Y (n5497) );
  OA21x2_ASAP7_75t_R   g5490( .A1 (n3989), .A2 (n5497), .B (n556), .Y (y2506) );
  AO21x1_ASAP7_75t_R   g5491( .A1 (n28), .A2 (x0), .B (n306), .Y (n5499) );
  AO21x1_ASAP7_75t_R   g5492( .A1 (x1), .A2 (n604), .B (n5499), .Y (y2507) );
  _const0_             g5493( .z (y2508) );
  AO32x1_ASAP7_75t_R   g5494( .A1 (y2079), .A2 (n108), .A3 (n155), .B1 (n763), .B2 (y232), .Y (y2509) );
  OA33x2_ASAP7_75t_R   g5495( .A1 (x0), .A2 (n671), .A3 (n403), .B1 (n22), .B2 (n628), .B3 (n421), .Y (y2510) );
  AO21x1_ASAP7_75t_R   g5496( .A1 (y2079), .A2 (n652), .B (n3189), .Y (y2511) );
  AND2x2_ASAP7_75t_R   g5497( .A (y1281), .B (n475), .Y (y2512) );
  AND2x2_ASAP7_75t_R   g5498( .A (n5145), .B (n3380), .Y (y2513) );
  OR3x1_ASAP7_75t_R    g5499( .A (x2), .B (x3), .C (x5), .Y (n5507) );
  AND2x2_ASAP7_75t_R   g5500( .A (y1474), .B (n5507), .Y (y2514) );
  AO21x1_ASAP7_75t_R   g5501( .A1 (n1163), .A2 (n3327), .B (n3055), .Y (y2515) );
  AND3x1_ASAP7_75t_R   g5502( .A (n776), .B (n740), .C (n12), .Y (n5510) );
  INVx1_ASAP7_75t_R    g5503( .A (n5510), .Y (y2516) );
  OR3x1_ASAP7_75t_R    g5504( .A (n1419), .B (n2070), .C (n143), .Y (y2517) );
  AO21x1_ASAP7_75t_R   g5505( .A1 (n310), .A2 (x3), .B (n3189), .Y (n5513) );
  OR3x1_ASAP7_75t_R    g5506( .A (n5513), .B (n3203), .C (x5), .Y (n5514) );
  INVx1_ASAP7_75t_R    g5507( .A (n5514), .Y (y2518) );
  NAND2x1_ASAP7_75t_R  g5508( .A (n12), .B (n391), .Y (n5516) );
  AO21x1_ASAP7_75t_R   g5509( .A1 (n5516), .A2 (y3293), .B (n959), .Y (y2519) );
  AND2x2_ASAP7_75t_R   g5510( .A (n23), .B (x3), .Y (n5518) );
  AO21x1_ASAP7_75t_R   g5511( .A1 (n4304), .A2 (x4), .B (n5518), .Y (y2520) );
  INVx1_ASAP7_75t_R    g5512( .A (n5173), .Y (n5520) );
  AND3x1_ASAP7_75t_R   g5513( .A (n5520), .B (n1572), .C (y2079), .Y (y2521) );
  INVx1_ASAP7_75t_R    g5514( .A (n638), .Y (n5522) );
  AND2x2_ASAP7_75t_R   g5515( .A (y1628), .B (n5522), .Y (y2522) );
  AND3x1_ASAP7_75t_R   g5516( .A (n968), .B (n219), .C (y2079), .Y (y2523) );
  AO21x1_ASAP7_75t_R   g5517( .A1 (n16), .A2 (n1373), .B (n1292), .Y (y2524) );
  AND3x1_ASAP7_75t_R   g5518( .A (y672), .B (n724), .C (y3377), .Y (y2525) );
  AND3x1_ASAP7_75t_R   g5519( .A (n4548), .B (n3459), .C (n401), .Y (y2526) );
  AO21x1_ASAP7_75t_R   g5520( .A1 (y2079), .A2 (n1342), .B (n337), .Y (y2527) );
  AO21x1_ASAP7_75t_R   g5521( .A1 (n3705), .A2 (n3918), .B (n45), .Y (n5529) );
  AND2x2_ASAP7_75t_R   g5522( .A (n5529), .B (n556), .Y (y2528) );
  NOR2x1_ASAP7_75t_R   g5523( .A (n756), .B (n290), .Y (n5531) );
  OR3x1_ASAP7_75t_R    g5524( .A (n5531), .B (n3279), .C (n628), .Y (y2529) );
  OR3x1_ASAP7_75t_R    g5525( .A (n1158), .B (n1775), .C (n2994), .Y (y2530) );
  AND2x2_ASAP7_75t_R   g5526( .A (n534), .B (y3852), .Y (n5534) );
  AO21x1_ASAP7_75t_R   g5527( .A1 (n497), .A2 (n5534), .B (n987), .Y (y2531) );
  NAND2x1_ASAP7_75t_R  g5528( .A (n558), .B (n3480), .Y (n5536) );
  AND2x2_ASAP7_75t_R   g5529( .A (n5536), .B (n1218), .Y (y2532) );
  AND2x2_ASAP7_75t_R   g5530( .A (n406), .B (n3089), .Y (y2533) );
  AND2x2_ASAP7_75t_R   g5531( .A (y3758), .B (x2), .Y (n5539) );
  AO21x1_ASAP7_75t_R   g5532( .A1 (n3618), .A2 (n3183), .B (n5539), .Y (y2534) );
  AND2x2_ASAP7_75t_R   g5533( .A (n415), .B (n4903), .Y (y2535) );
  AO21x1_ASAP7_75t_R   g5534( .A1 (n5520), .A2 (y2079), .B (n3316), .Y (y2536) );
  AO21x1_ASAP7_75t_R   g5535( .A1 (n137), .A2 (n72), .B (y2079), .Y (n5543) );
  INVx1_ASAP7_75t_R    g5536( .A (n5543), .Y (n5544) );
  OA33x2_ASAP7_75t_R   g5537( .A1 (x4), .A2 (n76), .A3 (n4575), .B1 (n22), .B2 (n5544), .B3 (n3963), .Y (y2537) );
  AND2x2_ASAP7_75t_R   g5538( .A (n868), .B (x0), .Y (y2538) );
  AO21x1_ASAP7_75t_R   g5539( .A1 (y2079), .A2 (x4), .B (n81), .Y (n5547) );
  AO21x1_ASAP7_75t_R   g5540( .A1 (n3860), .A2 (n5547), .B (n3135), .Y (y2539) );
  AND3x1_ASAP7_75t_R   g5541( .A (n369), .B (n290), .C (n343), .Y (y2540) );
  INVx1_ASAP7_75t_R    g5542( .A (n4155), .Y (n5550) );
  OA21x2_ASAP7_75t_R   g5543( .A1 (n5550), .A2 (x3), .B (n3882), .Y (y2541) );
  AND2x2_ASAP7_75t_R   g5544( .A (n4111), .B (y168), .Y (y2542) );
  AO21x1_ASAP7_75t_R   g5545( .A1 (x4), .A2 (n756), .B (y2466), .Y (n5553) );
  AO21x1_ASAP7_75t_R   g5546( .A1 (x3), .A2 (n4528), .B (n5553), .Y (n5554) );
  AND2x2_ASAP7_75t_R   g5547( .A (n5554), .B (n4241), .Y (y2543) );
  NAND2x1_ASAP7_75t_R  g5548( .A (x5), .B (n3989), .Y (y2648) );
  AND3x1_ASAP7_75t_R   g5549( .A (n337), .B (y2079), .C (n15), .Y (n5557) );
  INVx1_ASAP7_75t_R    g5550( .A (n5557), .Y (n5558) );
  AND2x2_ASAP7_75t_R   g5551( .A (y2648), .B (n5558), .Y (y2544) );
  AO21x1_ASAP7_75t_R   g5552( .A1 (n218), .A2 (n29), .B (n4459), .Y (y2545) );
  AO21x1_ASAP7_75t_R   g5553( .A1 (y2079), .A2 (n3792), .B (y1257), .Y (y2546) );
  INVx1_ASAP7_75t_R    g5554( .A (n1896), .Y (y2547) );
  AND2x2_ASAP7_75t_R   g5555( .A (n5279), .B (n2414), .Y (y2548) );
  AND2x2_ASAP7_75t_R   g5556( .A (n290), .B (y3852), .Y (n5564) );
  AO21x1_ASAP7_75t_R   g5557( .A1 (x4), .A2 (y2079), .B (n622), .Y (n5565) );
  AND2x2_ASAP7_75t_R   g5558( .A (n5564), .B (n5565), .Y (y2549) );
  AND2x2_ASAP7_75t_R   g5559( .A (n1863), .B (y2852), .Y (y2550) );
  AO21x1_ASAP7_75t_R   g5560( .A1 (y2079), .A2 (n22), .B (n76), .Y (n5568) );
  AND2x2_ASAP7_75t_R   g5561( .A (n4595), .B (n5568), .Y (n5569) );
  INVx1_ASAP7_75t_R    g5562( .A (n5569), .Y (y2551) );
  AND2x2_ASAP7_75t_R   g5563( .A (n4241), .B (n4276), .Y (y2552) );
  AO21x1_ASAP7_75t_R   g5564( .A1 (y2079), .A2 (x2), .B (n3847), .Y (y2553) );
  AO21x1_ASAP7_75t_R   g5565( .A1 (n3630), .A2 (x3), .B (n4925), .Y (y2554) );
  AO21x1_ASAP7_75t_R   g5566( .A1 (n388), .A2 (n3817), .B (x3), .Y (n5574) );
  AO21x1_ASAP7_75t_R   g5567( .A1 (n3567), .A2 (y2079), .B (n3338), .Y (n5575) );
  AND2x2_ASAP7_75t_R   g5568( .A (n5574), .B (n5575), .Y (y2555) );
  NOR2x1_ASAP7_75t_R   g5569( .A (n227), .B (n1541), .Y (y2556) );
  AO32x1_ASAP7_75t_R   g5570( .A1 (x1), .A2 (n746), .A3 (n1466), .B1 (n16), .B2 (n1889), .Y (y2557) );
  AND2x2_ASAP7_75t_R   g5571( .A (y1742), .B (n1851), .Y (y2558) );
  AO32x1_ASAP7_75t_R   g5572( .A1 (n1656), .A2 (x2), .A3 (n219), .B1 (n271), .B2 (n1657), .Y (y2559) );
  OA21x2_ASAP7_75t_R   g5573( .A1 (n2493), .A2 (n16), .B (n2503), .Y (y2560) );
  NAND2x1_ASAP7_75t_R  g5574( .A (n3256), .B (n4921), .Y (y2561) );
  AO21x1_ASAP7_75t_R   g5575( .A1 (y2079), .A2 (x3), .B (n3386), .Y (y2562) );
  AND3x1_ASAP7_75t_R   g5576( .A (n382), .B (n681), .C (y2079), .Y (y3305) );
  AO21x1_ASAP7_75t_R   g5577( .A1 (n22), .A2 (n421), .B (y3305), .Y (y2563) );
  AO21x1_ASAP7_75t_R   g5578( .A1 (y2079), .A2 (n310), .B (n3189), .Y (n5586) );
  NAND2x1_ASAP7_75t_R  g5579( .A (n671), .B (n299), .Y (n5587) );
  AND2x2_ASAP7_75t_R   g5580( .A (n5586), .B (n5587), .Y (y2564) );
  AO21x1_ASAP7_75t_R   g5581( .A1 (y2079), .A2 (n310), .B (n2718), .Y (n5589) );
  AND2x2_ASAP7_75t_R   g5582( .A (n5589), .B (n4907), .Y (y2565) );
  AO21x1_ASAP7_75t_R   g5583( .A1 (n753), .A2 (x0), .B (n701), .Y (y2566) );
  AO21x1_ASAP7_75t_R   g5584( .A1 (x0), .A2 (n4389), .B (n1860), .Y (y2567) );
  AO21x1_ASAP7_75t_R   g5585( .A1 (y2079), .A2 (n228), .B (n905), .Y (y2568) );
  AO21x1_ASAP7_75t_R   g5586( .A1 (y2079), .A2 (n3040), .B (n3189), .Y (y2569) );
  AO21x1_ASAP7_75t_R   g5587( .A1 (n4336), .A2 (y2079), .B (n2718), .Y (n5595) );
  AND2x2_ASAP7_75t_R   g5588( .A (n5595), .B (n4907), .Y (y2570) );
  AO21x1_ASAP7_75t_R   g5589( .A1 (y2079), .A2 (n4844), .B (n3751), .Y (y2571) );
  NOR2x1_ASAP7_75t_R   g5590( .A (n2756), .B (n1536), .Y (n5598) );
  AO21x1_ASAP7_75t_R   g5591( .A1 (n1676), .A2 (n17), .B (n5598), .Y (y2572) );
  AO21x1_ASAP7_75t_R   g5592( .A1 (n3121), .A2 (y2079), .B (n3386), .Y (y2573) );
  OA21x2_ASAP7_75t_R   g5593( .A1 (x2), .A2 (n5108), .B (n3209), .Y (y2574) );
  AO21x1_ASAP7_75t_R   g5594( .A1 (n3474), .A2 (n4375), .B (n4042), .Y (y2575) );
  OA21x2_ASAP7_75t_R   g5595( .A1 (n427), .A2 (n425), .B (n22), .Y (n5603) );
  AO21x1_ASAP7_75t_R   g5596( .A1 (n84), .A2 (n529), .B (n5603), .Y (y2576) );
  OA21x2_ASAP7_75t_R   g5597( .A1 (n2508), .A2 (n2146), .B (n2322), .Y (y2577) );
  AND3x1_ASAP7_75t_R   g5598( .A (n28), .B (n299), .C (n17), .Y (n5606) );
  NOR2x1_ASAP7_75t_R   g5599( .A (n3519), .B (n5606), .Y (y2579) );
  AND2x2_ASAP7_75t_R   g5600( .A (y2442), .B (n455), .Y (y2580) );
  INVx1_ASAP7_75t_R    g5601( .A (n3434), .Y (n5609) );
  AND3x1_ASAP7_75t_R   g5602( .A (n5609), .B (n1272), .C (n556), .Y (y2581) );
  AO21x1_ASAP7_75t_R   g5603( .A1 (n12), .A2 (y3293), .B (n297), .Y (n5611) );
  AO21x1_ASAP7_75t_R   g5604( .A1 (n5611), .A2 (n419), .B (n145), .Y (y2582) );
  NAND2x1_ASAP7_75t_R  g5605( .A (x4), .B (n4467), .Y (n5613) );
  AND3x1_ASAP7_75t_R   g5606( .A (n5613), .B (n2971), .C (n4638), .Y (y2583) );
  AND3x1_ASAP7_75t_R   g5607( .A (n382), .B (y3377), .C (x0), .Y (y2584) );
  OA211x2_ASAP7_75t_R  g5608( .A1 (n3116), .A2 (n3417), .B (n4559), .C (y3852), .Y (y2585) );
  OA21x2_ASAP7_75t_R   g5609( .A1 (n993), .A2 (n604), .B (n919), .Y (y2586) );
  AND2x2_ASAP7_75t_R   g5610( .A (n219), .B (n463), .Y (y2587) );
  AND2x2_ASAP7_75t_R   g5611( .A (n3445), .B (y2079), .Y (n5619) );
  AO21x1_ASAP7_75t_R   g5612( .A1 (n218), .A2 (n29), .B (n5619), .Y (y2588) );
  AO21x1_ASAP7_75t_R   g5613( .A1 (y2079), .A2 (n3989), .B (n4114), .Y (y2589) );
  AND2x2_ASAP7_75t_R   g5614( .A (y3377), .B (n330), .Y (y2590) );
  AO21x1_ASAP7_75t_R   g5615( .A1 (n93), .A2 (x0), .B (n787), .Y (y2591) );
  AND2x2_ASAP7_75t_R   g5616( .A (n189), .B (n406), .Y (y2592) );
  AO21x1_ASAP7_75t_R   g5617( .A1 (n164), .A2 (n173), .B (n262), .Y (y2593) );
  AND2x2_ASAP7_75t_R   g5618( .A (n4662), .B (n556), .Y (y2594) );
  OA21x2_ASAP7_75t_R   g5619( .A1 (n3502), .A2 (n552), .B (n2542), .Y (y2595) );
  AND3x1_ASAP7_75t_R   g5620( .A (n765), .B (n64), .C (n610), .Y (n5628) );
  NOR2x1_ASAP7_75t_R   g5621( .A (n1245), .B (n5628), .Y (y2596) );
  AO21x1_ASAP7_75t_R   g5622( .A1 (n3040), .A2 (y2079), .B (n347), .Y (n5630) );
  NOR2x1_ASAP7_75t_R   g5623( .A (y2079), .B (n4368), .Y (n5631) );
  AO21x1_ASAP7_75t_R   g5624( .A1 (n5056), .A2 (n5630), .B (n5631), .Y (y2597) );
  AND2x2_ASAP7_75t_R   g5625( .A (n360), .B (y2079), .Y (n5633) );
  OA21x2_ASAP7_75t_R   g5626( .A1 (n5633), .A2 (n3414), .B (n1620), .Y (y2598) );
  OR3x1_ASAP7_75t_R    g5627( .A (y1738), .B (n1501), .C (n2169), .Y (y2599) );
  OR3x1_ASAP7_75t_R    g5628( .A (n43), .B (n17), .C (x2), .Y (n5636) );
  INVx1_ASAP7_75t_R    g5629( .A (n5636), .Y (n5637) );
  OA21x2_ASAP7_75t_R   g5630( .A1 (n5637), .A2 (n143), .B (n2116), .Y (y2600) );
  AND2x2_ASAP7_75t_R   g5631( .A (y2632), .B (n4935), .Y (y2601) );
  INVx1_ASAP7_75t_R    g5632( .A (n349), .Y (n5640) );
  AO21x1_ASAP7_75t_R   g5633( .A1 (n319), .A2 (x4), .B (n426), .Y (n5641) );
  NAND2x1_ASAP7_75t_R  g5634( .A (n5640), .B (n5641), .Y (y2602) );
  INVx1_ASAP7_75t_R    g5635( .A (n3376), .Y (n5643) );
  AO21x1_ASAP7_75t_R   g5636( .A1 (n1062), .A2 (n5643), .B (n3847), .Y (y2603) );
  AND2x2_ASAP7_75t_R   g5637( .A (y3198), .B (n3884), .Y (y2604) );
  AO21x1_ASAP7_75t_R   g5638( .A1 (y2079), .A2 (n436), .B (n1150), .Y (y2605) );
  OR3x1_ASAP7_75t_R    g5639( .A (n914), .B (n403), .C (x5), .Y (n5647) );
  OA21x2_ASAP7_75t_R   g5640( .A1 (y2079), .A2 (n378), .B (n5647), .Y (y2606) );
  AO21x1_ASAP7_75t_R   g5641( .A1 (y2079), .A2 (n401), .B (n4349), .Y (y2608) );
  AO21x1_ASAP7_75t_R   g5642( .A1 (n12), .A2 (n534), .B (n1545), .Y (n5650) );
  INVx1_ASAP7_75t_R    g5643( .A (n5650), .Y (n5651) );
  AND2x2_ASAP7_75t_R   g5644( .A (n221), .B (y2079), .Y (n5652) );
  AO21x1_ASAP7_75t_R   g5645( .A1 (n455), .A2 (n5651), .B (n5652), .Y (y2609) );
  AO21x1_ASAP7_75t_R   g5646( .A1 (y2079), .A2 (x3), .B (n45), .Y (n5654) );
  AO21x1_ASAP7_75t_R   g5647( .A1 (x2), .A2 (n22), .B (n5654), .Y (y2610) );
  AND2x2_ASAP7_75t_R   g5648( .A (n2573), .B (n348), .Y (y2611) );
  AO21x1_ASAP7_75t_R   g5649( .A1 (n22), .A2 (n5176), .B (n4366), .Y (y2613) );
  AND2x2_ASAP7_75t_R   g5650( .A (n4755), .B (n4353), .Y (y2614) );
  NOR2x1_ASAP7_75t_R   g5651( .A (n12), .B (n1045), .Y (y2615) );
  NOR2x1_ASAP7_75t_R   g5652( .A (n2989), .B (n5438), .Y (y2616) );
  INVx1_ASAP7_75t_R    g5653( .A (n1917), .Y (n5661) );
  OA211x2_ASAP7_75t_R  g5654( .A1 (n5661), .A2 (n2843), .B (n3606), .C (n556), .Y (y2617) );
  AND3x1_ASAP7_75t_R   g5655( .A (n2116), .B (y3852), .C (n64), .Y (y2618) );
  AO21x1_ASAP7_75t_R   g5656( .A1 (n5181), .A2 (n2971), .B (n29), .Y (y2619) );
  NOR2x1_ASAP7_75t_R   g5657( .A (x5), .B (x2), .Y (n5665) );
  AO21x1_ASAP7_75t_R   g5658( .A1 (y2079), .A2 (n15), .B (x3), .Y (n5666) );
  NOR2x1_ASAP7_75t_R   g5659( .A (x4), .B (n5666), .Y (n5667) );
  AO21x1_ASAP7_75t_R   g5660( .A1 (n348), .A2 (n5665), .B (n5667), .Y (y2620) );
  AO21x1_ASAP7_75t_R   g5661( .A1 (n22), .A2 (n17), .B (n856), .Y (y2621) );
  OR4x2_ASAP7_75t_R    g5662( .A (n529), .B (n1032), .C (n2718), .D (x5), .Y (n5670) );
  AND2x2_ASAP7_75t_R   g5663( .A (y851), .B (n5670), .Y (y2622) );
  AO21x1_ASAP7_75t_R   g5664( .A1 (n63), .A2 (n3808), .B (n754), .Y (y2623) );
  INVx1_ASAP7_75t_R    g5665( .A (n489), .Y (n5673) );
  OA21x2_ASAP7_75t_R   g5666( .A1 (x1), .A2 (n5673), .B (n917), .Y (y2624) );
  OA21x2_ASAP7_75t_R   g5667( .A1 (n1278), .A2 (x2), .B (n3209), .Y (y2625) );
  AND2x2_ASAP7_75t_R   g5668( .A (n5516), .B (y3293), .Y (y2626) );
  AND3x1_ASAP7_75t_R   g5669( .A (n5296), .B (n3170), .C (n17), .Y (n5677) );
  INVx1_ASAP7_75t_R    g5670( .A (n5296), .Y (n5678) );
  INVx1_ASAP7_75t_R    g5671( .A (n3170), .Y (n5679) );
  OA21x2_ASAP7_75t_R   g5672( .A1 (n5678), .A2 (n5679), .B (x3), .Y (n5680) );
  OR2x4_ASAP7_75t_R    g5673( .A (n5677), .B (n5680), .Y (n5681) );
  AND2x2_ASAP7_75t_R   g5674( .A (n5681), .B (n4618), .Y (y2627) );
  OR3x1_ASAP7_75t_R    g5675( .A (n3443), .B (n15), .C (n337), .Y (n5683) );
  AND2x2_ASAP7_75t_R   g5676( .A (n5683), .B (n4129), .Y (y2628) );
  AO21x1_ASAP7_75t_R   g5677( .A1 (y3377), .A2 (n724), .B (x0), .Y (y2629) );
  INVx1_ASAP7_75t_R    g5678( .A (n1846), .Y (n5686) );
  AO21x1_ASAP7_75t_R   g5679( .A1 (n583), .A2 (n5686), .B (n1860), .Y (y2630) );
  AO21x1_ASAP7_75t_R   g5680( .A1 (n3469), .A2 (n3567), .B (n17), .Y (n5688) );
  INVx1_ASAP7_75t_R    g5681( .A (n5688), .Y (n5689) );
  INVx1_ASAP7_75t_R    g5682( .A (n3183), .Y (n5690) );
  AOI22x1_ASAP7_75t_R  g5683( .A1 (n5689), .A2 (n3183), .B1 (n5690), .B2 (n5688), .Y (y2631) );
  AND3x1_ASAP7_75t_R   g5684( .A (n17), .B (n22), .C (x2), .Y (n5692) );
  INVx1_ASAP7_75t_R    g5685( .A (n5692), .Y (n5693) );
  OA211x2_ASAP7_75t_R  g5686( .A1 (n4551), .A2 (y2079), .B (n3334), .C (n5693), .Y (y2633) );
  AND2x2_ASAP7_75t_R   g5687( .A (n2322), .B (n1562), .Y (y2634) );
  AND3x1_ASAP7_75t_R   g5688( .A (n28), .B (n137), .C (n72), .Y (n5696) );
  AO21x1_ASAP7_75t_R   g5689( .A1 (n218), .A2 (n29), .B (n5696), .Y (n5697) );
  NAND2x1_ASAP7_75t_R  g5690( .A (n316), .B (n5697), .Y (y2635) );
  AO32x1_ASAP7_75t_R   g5691( .A1 (y2079), .A2 (n401), .A3 (n72), .B1 (n1838), .B2 (n29), .Y (y2636) );
  INVx1_ASAP7_75t_R    g5692( .A (n5001), .Y (n5700) );
  AO21x1_ASAP7_75t_R   g5693( .A1 (x2), .A2 (y2079), .B (n290), .Y (n5701) );
  OA21x2_ASAP7_75t_R   g5694( .A1 (n5700), .A2 (n17), .B (n5701), .Y (y2637) );
  NAND2x1_ASAP7_75t_R  g5695( .A (n17), .B (n1635), .Y (n5703) );
  AO21x1_ASAP7_75t_R   g5696( .A1 (n17), .A2 (n1635), .B (n164), .Y (n5704) );
  AO32x1_ASAP7_75t_R   g5697( .A1 (n72), .A2 (n5703), .A3 (y435), .B1 (n221), .B2 (n5704), .Y (y2638) );
  AND3x1_ASAP7_75t_R   g5698( .A (n4662), .B (n3089), .C (n556), .Y (y2639) );
  AO21x1_ASAP7_75t_R   g5699( .A1 (n22), .A2 (x5), .B (n45), .Y (n5707) );
  AO21x1_ASAP7_75t_R   g5700( .A1 (y2079), .A2 (n3024), .B (n5707), .Y (y2640) );
  AND2x2_ASAP7_75t_R   g5701( .A (y3397), .B (n4695), .Y (y2641) );
  AO21x1_ASAP7_75t_R   g5702( .A1 (n1564), .A2 (n63), .B (n2347), .Y (y2642) );
  AO21x1_ASAP7_75t_R   g5703( .A1 (n299), .A2 (n17), .B (y1281), .Y (n5711) );
  AND2x2_ASAP7_75t_R   g5704( .A (n3212), .B (n5711), .Y (y2644) );
  AO21x1_ASAP7_75t_R   g5705( .A1 (n1240), .A2 (y2079), .B (n1708), .Y (y2645) );
  OR3x1_ASAP7_75t_R    g5706( .A (n3443), .B (n58), .C (n337), .Y (y2646) );
  AO21x1_ASAP7_75t_R   g5707( .A1 (n15), .A2 (n180), .B (n2165), .Y (y2647) );
  NAND2x1_ASAP7_75t_R  g5708( .A (n12), .B (n1407), .Y (n5716) );
  AND2x2_ASAP7_75t_R   g5709( .A (n5716), .B (n1246), .Y (y2649) );
  AO21x1_ASAP7_75t_R   g5710( .A1 (n455), .A2 (n3645), .B (n4403), .Y (n5718) );
  AND2x2_ASAP7_75t_R   g5711( .A (n5718), .B (n290), .Y (y2650) );
  NAND2x1_ASAP7_75t_R  g5712( .A (n227), .B (n740), .Y (n5720) );
  AND2x2_ASAP7_75t_R   g5713( .A (y535), .B (n5720), .Y (y2651) );
  OA22x2_ASAP7_75t_R   g5714( .A1 (n363), .A2 (n914), .B1 (n5072), .B2 (x4), .Y (y2652) );
  OR3x1_ASAP7_75t_R    g5715( .A (n495), .B (n798), .C (n791), .Y (y2653) );
  AO21x1_ASAP7_75t_R   g5716( .A1 (n1676), .A2 (y2079), .B (y2259), .Y (y2654) );
  AO21x1_ASAP7_75t_R   g5717( .A1 (n22), .A2 (n4304), .B (n4922), .Y (y2655) );
  AND2x2_ASAP7_75t_R   g5718( .A (y3852), .B (n93), .Y (y2656) );
  OR3x1_ASAP7_75t_R    g5719( .A (n378), .B (y2079), .C (n686), .Y (n5727) );
  OA21x2_ASAP7_75t_R   g5720( .A1 (n4061), .A2 (n330), .B (n5727), .Y (y2657) );
  AO21x1_ASAP7_75t_R   g5721( .A1 (n546), .A2 (n463), .B (n977), .Y (y2658) );
  AO21x1_ASAP7_75t_R   g5722( .A1 (n22), .A2 (x5), .B (x3), .Y (n5730) );
  AND2x2_ASAP7_75t_R   g5723( .A (n3645), .B (n5730), .Y (y2660) );
  AO21x1_ASAP7_75t_R   g5724( .A1 (x1), .A2 (x3), .B (n12), .Y (n5732) );
  INVx1_ASAP7_75t_R    g5725( .A (n5732), .Y (n5733) );
  INVx1_ASAP7_75t_R    g5726( .A (n874), .Y (n5734) );
  NOR2x1_ASAP7_75t_R   g5727( .A (n12), .B (n4253), .Y (n5735) );
  INVx1_ASAP7_75t_R    g5728( .A (n5735), .Y (n5736) );
  OA211x2_ASAP7_75t_R  g5729( .A1 (n5733), .A2 (n5734), .B (n5736), .C (n84), .Y (y2661) );
  AO21x1_ASAP7_75t_R   g5730( .A1 (x3), .A2 (x5), .B (x2), .Y (n5738) );
  INVx1_ASAP7_75t_R    g5731( .A (n5738), .Y (n5739) );
  AO21x1_ASAP7_75t_R   g5732( .A1 (n4089), .A2 (n1572), .B (x4), .Y (n5740) );
  OA21x2_ASAP7_75t_R   g5733( .A1 (n5739), .A2 (n370), .B (n5740), .Y (y2662) );
  AND2x2_ASAP7_75t_R   g5734( .A (n4469), .B (y1359), .Y (y2663) );
  AND3x1_ASAP7_75t_R   g5735( .A (y1903), .B (n656), .C (n401), .Y (y2664) );
  INVx1_ASAP7_75t_R    g5736( .A (n868), .Y (n5744) );
  NOR2x1_ASAP7_75t_R   g5737( .A (n2738), .B (n2742), .Y (y2916) );
  AO21x1_ASAP7_75t_R   g5738( .A1 (n5744), .A2 (n12), .B (y2916), .Y (y2665) );
  AND2x2_ASAP7_75t_R   g5739( .A (y1474), .B (n3526), .Y (y2666) );
  AND2x2_ASAP7_75t_R   g5740( .A (y1903), .B (n3166), .Y (y2667) );
  AO21x1_ASAP7_75t_R   g5741( .A1 (n455), .A2 (y3852), .B (n3423), .Y (y2668) );
  AND3x1_ASAP7_75t_R   g5742( .A (n3705), .B (n5507), .C (n556), .Y (y2669) );
  NAND2x1_ASAP7_75t_R  g5743( .A (n388), .B (n3134), .Y (y2670) );
  INVx1_ASAP7_75t_R    g5744( .A (n4033), .Y (n5752) );
  OR3x1_ASAP7_75t_R    g5745( .A (n29), .B (n5752), .C (n45), .Y (y2671) );
  AO21x1_ASAP7_75t_R   g5746( .A1 (y9), .A2 (n312), .B (x4), .Y (n5754) );
  AND2x2_ASAP7_75t_R   g5747( .A (n5754), .B (n556), .Y (y2672) );
  OR3x1_ASAP7_75t_R    g5748( .A (x2), .B (x4), .C (x5), .Y (n5756) );
  AND3x1_ASAP7_75t_R   g5749( .A (n5442), .B (n369), .C (n5756), .Y (y2673) );
  AO21x1_ASAP7_75t_R   g5750( .A1 (n746), .A2 (x3), .B (n747), .Y (n5758) );
  AO21x1_ASAP7_75t_R   g5751( .A1 (n84), .A2 (n15), .B (n611), .Y (n5759) );
  AOI21x1_ASAP7_75t_R  g5752( .A1 (n5758), .A2 (n5759), .B (n2423), .Y (y2674) );
  AO32x1_ASAP7_75t_R   g5753( .A1 (n672), .A2 (n660), .A3 (x0), .B1 (y2079), .B2 (n3792), .Y (y2675) );
  AND3x1_ASAP7_75t_R   g5754( .A (n72), .B (n137), .C (n3029), .Y (y2676) );
  OR3x1_ASAP7_75t_R    g5755( .A (x1), .B (x0), .C (x3), .Y (n5763) );
  INVx1_ASAP7_75t_R    g5756( .A (n5763), .Y (n5764) );
  AO21x1_ASAP7_75t_R   g5757( .A1 (n5764), .A2 (n15), .B (y319), .Y (y2677) );
  NOR2x1_ASAP7_75t_R   g5758( .A (x1), .B (n2140), .Y (n5766) );
  INVx1_ASAP7_75t_R    g5759( .A (n5766), .Y (n5767) );
  AO21x1_ASAP7_75t_R   g5760( .A1 (n776), .A2 (n841), .B (x0), .Y (n5768) );
  AND2x2_ASAP7_75t_R   g5761( .A (n5767), .B (n5768), .Y (y2678) );
  AND2x2_ASAP7_75t_R   g5762( .A (n556), .B (n4099), .Y (n5770) );
  AO21x1_ASAP7_75t_R   g5763( .A1 (n352), .A2 (n5770), .B (n4922), .Y (y2679) );
  AND2x2_ASAP7_75t_R   g5764( .A (y1903), .B (n4249), .Y (y2680) );
  AO21x1_ASAP7_75t_R   g5765( .A1 (n388), .A2 (n28), .B (n137), .Y (n5773) );
  AND3x1_ASAP7_75t_R   g5766( .A (n5773), .B (n3119), .C (n5756), .Y (y2681) );
  AO21x1_ASAP7_75t_R   g5767( .A1 (n312), .A2 (n497), .B (x0), .Y (n5775) );
  NOR2x1_ASAP7_75t_R   g5768( .A (x2), .B (n5775), .Y (n5776) );
  AND2x2_ASAP7_75t_R   g5769( .A (n1066), .B (n800), .Y (n5777) );
  OR3x1_ASAP7_75t_R    g5770( .A (n5776), .B (n5777), .C (y2196), .Y (y2682) );
  AO21x1_ASAP7_75t_R   g5771( .A1 (n334), .A2 (y2079), .B (n337), .Y (n5779) );
  AND2x2_ASAP7_75t_R   g5772( .A (n5779), .B (n3979), .Y (y2683) );
  AO21x1_ASAP7_75t_R   g5773( .A1 (n556), .A2 (n5090), .B (n3263), .Y (y2684) );
  AND3x1_ASAP7_75t_R   g5774( .A (n3966), .B (n858), .C (n497), .Y (y2685) );
  AO21x1_ASAP7_75t_R   g5775( .A1 (y2079), .A2 (x2), .B (n3025), .Y (y2872) );
  AND2x2_ASAP7_75t_R   g5776( .A (y2872), .B (n4171), .Y (y2686) );
  AND3x1_ASAP7_75t_R   g5777( .A (n4329), .B (n1838), .C (n556), .Y (y2687) );
  OA21x2_ASAP7_75t_R   g5778( .A1 (x3), .A2 (n308), .B (n3882), .Y (y2688) );
  AO21x1_ASAP7_75t_R   g5779( .A1 (n178), .A2 (x0), .B (n787), .Y (y2689) );
  AO21x1_ASAP7_75t_R   g5780( .A1 (n527), .A2 (n352), .B (n957), .Y (y2690) );
  AND2x2_ASAP7_75t_R   g5781( .A (n1191), .B (n1272), .Y (y2691) );
  AND2x2_ASAP7_75t_R   g5782( .A (n2577), .B (n2726), .Y (n5790) );
  AND3x1_ASAP7_75t_R   g5783( .A (n5790), .B (n64), .C (n63), .Y (y2692) );
  AO21x1_ASAP7_75t_R   g5784( .A1 (n17), .A2 (n341), .B (n3234), .Y (y2693) );
  AO21x1_ASAP7_75t_R   g5785( .A1 (y2079), .A2 (n3448), .B (n4878), .Y (y2694) );
  AO21x1_ASAP7_75t_R   g5786( .A1 (n989), .A2 (x2), .B (n1644), .Y (y2695) );
  AND2x2_ASAP7_75t_R   g5787( .A (n4111), .B (n4933), .Y (y2696) );
  AND2x2_ASAP7_75t_R   g5788( .A (n4933), .B (n645), .Y (y2697) );
  OA21x2_ASAP7_75t_R   g5789( .A1 (n2647), .A2 (n747), .B (n2465), .Y (y2698) );
  AO21x1_ASAP7_75t_R   g5790( .A1 (n22), .A2 (n583), .B (n1817), .Y (n5798) );
  AO32x1_ASAP7_75t_R   g5791( .A1 (x3), .A2 (n299), .A3 (y2079), .B1 (n17), .B2 (n5798), .Y (y2699) );
  AO21x1_ASAP7_75t_R   g5792( .A1 (n28), .A2 (n388), .B (n17), .Y (n5800) );
  AO21x1_ASAP7_75t_R   g5793( .A1 (y2079), .A2 (x4), .B (x3), .Y (n5801) );
  OR3x1_ASAP7_75t_R    g5794( .A (n29), .B (n5801), .C (n12), .Y (n5802) );
  NAND2x1_ASAP7_75t_R  g5795( .A (n5800), .B (n5802), .Y (y2700) );
  AND2x2_ASAP7_75t_R   g5796( .A (y2727), .B (n672), .Y (y2701) );
  AO21x1_ASAP7_75t_R   g5797( .A1 (n5345), .A2 (y2079), .B (n638), .Y (y2702) );
  AO21x1_ASAP7_75t_R   g5798( .A1 (n836), .A2 (y3852), .B (n713), .Y (y2703) );
  NOR2x1_ASAP7_75t_R   g5799( .A (n1927), .B (n3390), .Y (y2704) );
  INVx1_ASAP7_75t_R    g5800( .A (n4528), .Y (n5808) );
  AND3x1_ASAP7_75t_R   g5801( .A (n369), .B (n290), .C (x2), .Y (n5809) );
  AO21x1_ASAP7_75t_R   g5802( .A1 (n678), .A2 (n5808), .B (n5809), .Y (y2705) );
  AO21x1_ASAP7_75t_R   g5803( .A1 (x3), .A2 (n22), .B (n4972), .Y (n5811) );
  INVx1_ASAP7_75t_R    g5804( .A (n5811), .Y (n5812) );
  OA21x2_ASAP7_75t_R   g5805( .A1 (n5812), .A2 (n4486), .B (n3030), .Y (y2706) );
  AND2x2_ASAP7_75t_R   g5806( .A (n899), .B (y2079), .Y (y2707) );
  AO21x1_ASAP7_75t_R   g5807( .A1 (y2079), .A2 (x0), .B (n4250), .Y (y2708) );
  OR3x1_ASAP7_75t_R    g5808( .A (n999), .B (n12), .C (x5), .Y (n5816) );
  AND2x2_ASAP7_75t_R   g5809( .A (n5816), .B (y136), .Y (y2709) );
  AO21x1_ASAP7_75t_R   g5810( .A1 (n1564), .A2 (n63), .B (n2440), .Y (y2710) );
  INVx1_ASAP7_75t_R    g5811( .A (n4487), .Y (n5819) );
  AO21x1_ASAP7_75t_R   g5812( .A1 (n5819), .A2 (y2079), .B (n4514), .Y (y2711) );
  OA21x2_ASAP7_75t_R   g5813( .A1 (n2647), .A2 (n1255), .B (n2414), .Y (y2712) );
  AND2x2_ASAP7_75t_R   g5814( .A (n3109), .B (y3176), .Y (y2713) );
  AND2x2_ASAP7_75t_R   g5815( .A (n4083), .B (n219), .Y (y2714) );
  AND3x1_ASAP7_75t_R   g5816( .A (n72), .B (n4495), .C (y2079), .Y (y3883) );
  INVx1_ASAP7_75t_R    g5817( .A (y3883), .Y (n5825) );
  AND2x2_ASAP7_75t_R   g5818( .A (n5825), .B (y3171), .Y (y2715) );
  AND3x1_ASAP7_75t_R   g5819( .A (x4), .B (x3), .C (x5), .Y (n5827) );
  INVx1_ASAP7_75t_R    g5820( .A (n5827), .Y (n5828) );
  AND3x1_ASAP7_75t_R   g5821( .A (n5493), .B (n5828), .C (n652), .Y (y2717) );
  NAND2x1_ASAP7_75t_R  g5822( .A (x5), .B (n5465), .Y (n5830) );
  AND2x2_ASAP7_75t_R   g5823( .A (n5830), .B (n4789), .Y (y2718) );
  NAND2x1_ASAP7_75t_R  g5824( .A (n16), .B (n1047), .Y (n5832) );
  AO21x1_ASAP7_75t_R   g5825( .A1 (n388), .A2 (n961), .B (x0), .Y (n5833) );
  OA21x2_ASAP7_75t_R   g5826( .A1 (y3758), .A2 (n5832), .B (n5833), .Y (y2719) );
  AO21x1_ASAP7_75t_R   g5827( .A1 (n421), .A2 (n3028), .B (n3630), .Y (y2720) );
  AO21x1_ASAP7_75t_R   g5828( .A1 (n4564), .A2 (x3), .B (n3657), .Y (y2721) );
  AO21x1_ASAP7_75t_R   g5829( .A1 (y1693), .A2 (x2), .B (n3333), .Y (y2722) );
  AO21x1_ASAP7_75t_R   g5830( .A1 (n1775), .A2 (x3), .B (n3386), .Y (y2724) );
  AND2x2_ASAP7_75t_R   g5831( .A (n352), .B (y3852), .Y (n5839) );
  INVx1_ASAP7_75t_R    g5832( .A (n5839), .Y (n5840) );
  AO21x1_ASAP7_75t_R   g5833( .A1 (n352), .A2 (n103), .B (n128), .Y (n5841) );
  XOR2x2_ASAP7_75t_R   g5834( .A (n5840), .B (n5841), .Y (y2725) );
  NAND2x1_ASAP7_75t_R  g5835( .A (x5), .B (n334), .Y (n5843) );
  OA21x2_ASAP7_75t_R   g5836( .A1 (n4920), .A2 (n3376), .B (n5843), .Y (y2726) );
  AO21x1_ASAP7_75t_R   g5837( .A1 (n1640), .A2 (n64), .B (x0), .Y (y2728) );
  OR3x1_ASAP7_75t_R    g5838( .A (n296), .B (n297), .C (y2498), .Y (y2729) );
  AO21x1_ASAP7_75t_R   g5839( .A1 (n29), .A2 (n77), .B (n3132), .Y (y2730) );
  OA21x2_ASAP7_75t_R   g5840( .A1 (n2610), .A2 (n495), .B (n1624), .Y (y2731) );
  AO21x1_ASAP7_75t_R   g5841( .A1 (y2079), .A2 (n3804), .B (n4460), .Y (y2732) );
  OA21x2_ASAP7_75t_R   g5842( .A1 (n4494), .A2 (n5314), .B (n3302), .Y (y2733) );
  AO21x1_ASAP7_75t_R   g5843( .A1 (n740), .A2 (n337), .B (n3443), .Y (y2734) );
  AND3x1_ASAP7_75t_R   g5844( .A (n4083), .B (n219), .C (n556), .Y (y2735) );
  AND3x1_ASAP7_75t_R   g5845( .A (n84), .B (n125), .C (x4), .Y (n5853) );
  INVx1_ASAP7_75t_R    g5846( .A (n5853), .Y (n5854) );
  NOR2x1_ASAP7_75t_R   g5847( .A (x3), .B (n3480), .Y (n5855) );
  AO21x1_ASAP7_75t_R   g5848( .A1 (n5854), .A2 (n4048), .B (n5855), .Y (y2736) );
  NAND2x1_ASAP7_75t_R  g5849( .A (x5), .B (n2989), .Y (n5857) );
  INVx1_ASAP7_75t_R    g5850( .A (n5857), .Y (n5858) );
  NOR2x1_ASAP7_75t_R   g5851( .A (x5), .B (n2989), .Y (n5859) );
  OR3x1_ASAP7_75t_R    g5852( .A (n5858), .B (n5859), .C (n45), .Y (y2738) );
  AND2x2_ASAP7_75t_R   g5853( .A (y2197), .B (n5094), .Y (y2741) );
  NAND2x1_ASAP7_75t_R  g5854( .A (n5116), .B (n285), .Y (n5862) );
  OA21x2_ASAP7_75t_R   g5855( .A1 (n3310), .A2 (n5862), .B (n4643), .Y (y2742) );
  AO21x1_ASAP7_75t_R   g5856( .A1 (n628), .A2 (n1851), .B (n337), .Y (y2743) );
  NOR2x1_ASAP7_75t_R   g5857( .A (n4486), .B (n4644), .Y (y2744) );
  AO21x1_ASAP7_75t_R   g5858( .A1 (n4618), .A2 (n4619), .B (n4047), .Y (y2745) );
  NAND2x1_ASAP7_75t_R  g5859( .A (y2079), .B (n5116), .Y (n5867) );
  INVx1_ASAP7_75t_R    g5860( .A (n5867), .Y (n5868) );
  AO21x1_ASAP7_75t_R   g5861( .A1 (n15), .A2 (y2079), .B (x3), .Y (n5869) );
  NOR2x1_ASAP7_75t_R   g5862( .A (x4), .B (n5869), .Y (n5870) );
  AO21x1_ASAP7_75t_R   g5863( .A1 (n348), .A2 (n5868), .B (n5870), .Y (y2746) );
  OA21x2_ASAP7_75t_R   g5864( .A1 (n3637), .A2 (n3918), .B (n406), .Y (y2747) );
  OA21x2_ASAP7_75t_R   g5865( .A1 (x0), .A2 (n1190), .B (n1001), .Y (y2748) );
  AO21x1_ASAP7_75t_R   g5866( .A1 (n137), .A2 (y2079), .B (n337), .Y (y2749) );
  AND2x2_ASAP7_75t_R   g5867( .A (n5103), .B (n406), .Y (y2750) );
  NOR2x1_ASAP7_75t_R   g5868( .A (x5), .B (n3143), .Y (n5876) );
  INVx1_ASAP7_75t_R    g5869( .A (n5876), .Y (n5877) );
  AND2x2_ASAP7_75t_R   g5870( .A (n5877), .B (n3919), .Y (y2751) );
  AO21x1_ASAP7_75t_R   g5871( .A1 (n660), .A2 (n137), .B (y2079), .Y (n5879) );
  AND2x2_ASAP7_75t_R   g5872( .A (n5879), .B (n3491), .Y (y2752) );
  AND2x2_ASAP7_75t_R   g5873( .A (n4548), .B (n72), .Y (y2753) );
  AO21x1_ASAP7_75t_R   g5874( .A1 (n3338), .A2 (n299), .B (n3417), .Y (y2754) );
  AO32x1_ASAP7_75t_R   g5875( .A1 (n299), .A2 (n1166), .A3 (x5), .B1 (n501), .B2 (n913), .Y (y2755) );
  AND2x2_ASAP7_75t_R   g5876( .A (n5085), .B (x3), .Y (n5884) );
  OA21x2_ASAP7_75t_R   g5877( .A1 (n5884), .A2 (n4981), .B (n4419), .Y (y2756) );
  AND3x1_ASAP7_75t_R   g5878( .A (n363), .B (n17), .C (n22), .Y (n5886) );
  NOR2x1_ASAP7_75t_R   g5879( .A (n5886), .B (n4486), .Y (y2757) );
  AO21x1_ASAP7_75t_R   g5880( .A1 (n378), .A2 (x0), .B (n2051), .Y (y2758) );
  NAND2x1_ASAP7_75t_R  g5881( .A (x3), .B (n3780), .Y (n5889) );
  AO21x1_ASAP7_75t_R   g5882( .A1 (n5889), .A2 (n137), .B (n418), .Y (y3100) );
  AND2x2_ASAP7_75t_R   g5883( .A (y3100), .B (n4632), .Y (y2759) );
  OR3x1_ASAP7_75t_R    g5884( .A (n139), .B (y2079), .C (n22), .Y (n5892) );
  AND2x2_ASAP7_75t_R   g5885( .A (n5892), .B (n343), .Y (n5893) );
  INVx1_ASAP7_75t_R    g5886( .A (n4065), .Y (n5894) );
  AOI21x1_ASAP7_75t_R  g5887( .A1 (n17), .A2 (n5893), .B (n5894), .Y (y2760) );
  OA21x2_ASAP7_75t_R   g5888( .A1 (n529), .A2 (n661), .B (n4508), .Y (y2761) );
  OR3x1_ASAP7_75t_R    g5889( .A (n5425), .B (n1029), .C (n529), .Y (y2762) );
  AND3x1_ASAP7_75t_R   g5890( .A (n413), .B (n348), .C (y2079), .Y (y2763) );
  AND3x1_ASAP7_75t_R   g5891( .A (n534), .B (n299), .C (y2079), .Y (y2764) );
  AO21x1_ASAP7_75t_R   g5892( .A1 (n1208), .A2 (y3293), .B (n4047), .Y (y2765) );
  NOR2x1_ASAP7_75t_R   g5893( .A (n3447), .B (n3677), .Y (y2766) );
  AND2x2_ASAP7_75t_R   g5894( .A (n1213), .B (x0), .Y (y2767) );
  AO21x1_ASAP7_75t_R   g5895( .A1 (n244), .A2 (n746), .B (x1), .Y (n5903) );
  INVx1_ASAP7_75t_R    g5896( .A (n5903), .Y (n5904) );
  INVx1_ASAP7_75t_R    g5897( .A (n692), .Y (n5905) );
  OA21x2_ASAP7_75t_R   g5898( .A1 (n5905), .A2 (n2070), .B (x1), .Y (n5906) );
  AO21x1_ASAP7_75t_R   g5899( .A1 (n5904), .A2 (y2079), .B (n5906), .Y (y2768) );
  AO21x1_ASAP7_75t_R   g5900( .A1 (n228), .A2 (n529), .B (n905), .Y (y2769) );
  AND2x2_ASAP7_75t_R   g5901( .A (n4109), .B (n556), .Y (y2772) );
  OR3x1_ASAP7_75t_R    g5902( .A (n81), .B (y2079), .C (n22), .Y (n5910) );
  OA21x2_ASAP7_75t_R   g5903( .A1 (n3859), .A2 (n3282), .B (n5910), .Y (y2773) );
  AND3x1_ASAP7_75t_R   g5904( .A (n818), .B (n819), .C (n895), .Y (y2774) );
  NAND2x1_ASAP7_75t_R  g5905( .A (n614), .B (n3077), .Y (y2775) );
  OA21x2_ASAP7_75t_R   g5906( .A1 (n999), .A2 (n1247), .B (n3380), .Y (y2776) );
  AO21x1_ASAP7_75t_R   g5907( .A1 (n5422), .A2 (y2079), .B (n300), .Y (y2777) );
  NAND2x1_ASAP7_75t_R  g5908( .A (x4), .B (n3866), .Y (n5916) );
  AND2x2_ASAP7_75t_R   g5909( .A (n5916), .B (n4109), .Y (y2779) );
  OR3x1_ASAP7_75t_R    g5910( .A (n3637), .B (n3918), .C (n337), .Y (n5918) );
  AND2x2_ASAP7_75t_R   g5911( .A (n5918), .B (y1693), .Y (y2780) );
  AND2x2_ASAP7_75t_R   g5912( .A (n656), .B (y2727), .Y (y2781) );
  AO21x1_ASAP7_75t_R   g5913( .A1 (n1432), .A2 (n22), .B (n349), .Y (y2782) );
  AO21x1_ASAP7_75t_R   g5914( .A1 (n3191), .A2 (n474), .B (n3129), .Y (y2783) );
  AO32x1_ASAP7_75t_R   g5915( .A1 (n388), .A2 (n3763), .A3 (n369), .B1 (x2), .B2 (y3758), .Y (y2784) );
  AOI21x1_ASAP7_75t_R  g5916( .A1 (n1838), .A2 (n1688), .B (n1653), .Y (y2785) );
  NOR2x1_ASAP7_75t_R   g5917( .A (n4586), .B (n1927), .Y (y2786) );
  AND3x1_ASAP7_75t_R   g5918( .A (n299), .B (n17), .C (x5), .Y (n5926) );
  AO21x1_ASAP7_75t_R   g5919( .A1 (n5493), .A2 (y1281), .B (n5926), .Y (y2788) );
  AO21x1_ASAP7_75t_R   g5920( .A1 (n15), .A2 (y2079), .B (n17), .Y (n5928) );
  INVx1_ASAP7_75t_R    g5921( .A (n5928), .Y (n5929) );
  AOI221x1_ASAP7_75t_R g5922( .A1 (n3025), .A2 (n3023), .B1 (n4695), .B2 (n5929), .C (n518), .Y (y2789) );
  AO21x1_ASAP7_75t_R   g5923( .A1 (n3000), .A2 (y2079), .B (n3338), .Y (n5931) );
  AO21x1_ASAP7_75t_R   g5924( .A1 (n28), .A2 (n740), .B (x3), .Y (n5932) );
  AND2x2_ASAP7_75t_R   g5925( .A (n5931), .B (n5932), .Y (y2790) );
  OA21x2_ASAP7_75t_R   g5926( .A1 (n3268), .A2 (n3269), .B (n556), .Y (y2791) );
  OA21x2_ASAP7_75t_R   g5927( .A1 (n1269), .A2 (n1457), .B (n844), .Y (y2792) );
  AO21x1_ASAP7_75t_R   g5928( .A1 (n22), .A2 (n1066), .B (n1907), .Y (y2793) );
  AND2x2_ASAP7_75t_R   g5929( .A (y2737), .B (n4732), .Y (y2794) );
  AND2x2_ASAP7_75t_R   g5930( .A (n3278), .B (n4439), .Y (y2795) );
  OR3x1_ASAP7_75t_R    g5931( .A (y2466), .B (n17), .C (n15), .Y (n5939) );
  AND3x1_ASAP7_75t_R   g5932( .A (n4329), .B (n5939), .C (n556), .Y (y2796) );
  AO21x1_ASAP7_75t_R   g5933( .A1 (n968), .A2 (n1077), .B (y2079), .Y (n5941) );
  OR3x1_ASAP7_75t_R    g5934( .A (n537), .B (x5), .C (x1), .Y (n5942) );
  AND2x2_ASAP7_75t_R   g5935( .A (n5941), .B (n5942), .Y (y2797) );
  AO21x1_ASAP7_75t_R   g5936( .A1 (n2971), .A2 (n4638), .B (n3316), .Y (y2798) );
  AO21x1_ASAP7_75t_R   g5937( .A1 (n16), .A2 (n812), .B (y2538), .Y (y2799) );
  AO21x1_ASAP7_75t_R   g5938( .A1 (n22), .A2 (n3191), .B (n3073), .Y (y2800) );
  AO21x1_ASAP7_75t_R   g5939( .A1 (n22), .A2 (n3192), .B (n3415), .Y (y2801) );
  AND3x1_ASAP7_75t_R   g5940( .A (n5939), .B (n556), .C (n3526), .Y (y2802) );
  AO21x1_ASAP7_75t_R   g5941( .A1 (n112), .A2 (n113), .B (n192), .Y (y2803) );
  AND2x2_ASAP7_75t_R   g5942( .A (n3327), .B (n4305), .Y (y2804) );
  INVx1_ASAP7_75t_R    g5943( .A (n247), .Y (n5951) );
  AO21x1_ASAP7_75t_R   g5944( .A1 (n17), .A2 (x0), .B (n1253), .Y (n5952) );
  AO32x1_ASAP7_75t_R   g5945( .A1 (n125), .A2 (n5951), .A3 (x1), .B1 (n1301), .B2 (n5952), .Y (y2805) );
  AND2x2_ASAP7_75t_R   g5946( .A (n3446), .B (n5303), .Y (y2806) );
  AND2x2_ASAP7_75t_R   g5947( .A (y3132), .B (x0), .Y (y2807) );
  OR3x1_ASAP7_75t_R    g5948( .A (n1261), .B (n1262), .C (n17), .Y (n5956) );
  NAND2x1_ASAP7_75t_R  g5949( .A (n797), .B (n5956), .Y (n5957) );
  AO21x1_ASAP7_75t_R   g5950( .A1 (n1613), .A2 (n17), .B (n5957), .Y (y2808) );
  AO21x1_ASAP7_75t_R   g5951( .A1 (n12), .A2 (y2079), .B (n3189), .Y (y2809) );
  NOR2x1_ASAP7_75t_R   g5952( .A (n392), .B (n959), .Y (y2810) );
  OA21x2_ASAP7_75t_R   g5953( .A1 (n3899), .A2 (n4459), .B (n1572), .Y (y2811) );
  OA21x2_ASAP7_75t_R   g5954( .A1 (n4139), .A2 (n1399), .B (n419), .Y (y2812) );
  INVx1_ASAP7_75t_R    g5955( .A (n3192), .Y (n5963) );
  AO21x1_ASAP7_75t_R   g5956( .A1 (n5963), .A2 (n84), .B (x4), .Y (n5964) );
  OA21x2_ASAP7_75t_R   g5957( .A1 (n22), .A2 (n3193), .B (n5964), .Y (y2814) );
  OR3x1_ASAP7_75t_R    g5958( .A (n581), .B (n1093), .C (n563), .Y (y2816) );
  OR3x1_ASAP7_75t_R    g5959( .A (n1158), .B (n4527), .C (n297), .Y (y3754) );
  INVx1_ASAP7_75t_R    g5960( .A (y3754), .Y (n5968) );
  NOR2x1_ASAP7_75t_R   g5961( .A (n15), .B (n5968), .Y (n5969) );
  AO21x1_ASAP7_75t_R   g5962( .A1 (n15), .A2 (n5968), .B (n5969), .Y (y2817) );
  OA21x2_ASAP7_75t_R   g5963( .A1 (n5544), .A2 (n5619), .B (n2998), .Y (y2818) );
  AND3x1_ASAP7_75t_R   g5964( .A (n4416), .B (n3780), .C (n17), .Y (n5972) );
  AO21x1_ASAP7_75t_R   g5965( .A1 (n391), .A2 (n4417), .B (n5972), .Y (y2819) );
  AO21x1_ASAP7_75t_R   g5966( .A1 (n1269), .A2 (n348), .B (n4868), .Y (y2820) );
  AND2x2_ASAP7_75t_R   g5967( .A (y1110), .B (n1894), .Y (y2821) );
  AND2x2_ASAP7_75t_R   g5968( .A (n534), .B (n299), .Y (n5976) );
  AO21x1_ASAP7_75t_R   g5969( .A1 (n466), .A2 (n363), .B (n5976), .Y (y2822) );
  AND3x1_ASAP7_75t_R   g5970( .A (n455), .B (n757), .C (n3469), .Y (n5978) );
  OA21x2_ASAP7_75t_R   g5971( .A1 (n5978), .A2 (n17), .B (n3181), .Y (y2823) );
  AO21x1_ASAP7_75t_R   g5972( .A1 (n17), .A2 (x1), .B (x2), .Y (n5980) );
  AO21x1_ASAP7_75t_R   g5973( .A1 (n189), .A2 (n16), .B (n5980), .Y (n5981) );
  OA21x2_ASAP7_75t_R   g5974( .A1 (n2565), .A2 (n202), .B (n5981), .Y (y2824) );
  AND2x2_ASAP7_75t_R   g5975( .A (y2450), .B (n453), .Y (y2825) );
  AND2x2_ASAP7_75t_R   g5976( .A (y3377), .B (x0), .Y (y2827) );
  AND3x1_ASAP7_75t_R   g5977( .A (n14), .B (n108), .C (y2079), .Y (n5985) );
  NOR2x1_ASAP7_75t_R   g5978( .A (n481), .B (n5985), .Y (y2828) );
  NAND2x1_ASAP7_75t_R  g5979( .A (n22), .B (n354), .Y (n5987) );
  AND3x1_ASAP7_75t_R   g5980( .A (n5987), .B (y1281), .C (n290), .Y (y2829) );
  AO21x1_ASAP7_75t_R   g5981( .A1 (n4321), .A2 (n3119), .B (n3427), .Y (y2830) );
  AO21x1_ASAP7_75t_R   g5982( .A1 (n856), .A2 (n17), .B (n22), .Y (n5990) );
  AND3x1_ASAP7_75t_R   g5983( .A (n4031), .B (n5990), .C (n3023), .Y (y2831) );
  AO21x1_ASAP7_75t_R   g5984( .A1 (n5250), .A2 (x2), .B (n45), .Y (y2833) );
  NAND2x1_ASAP7_75t_R  g5985( .A (x4), .B (n5177), .Y (n5993) );
  AND3x1_ASAP7_75t_R   g5986( .A (n671), .B (n22), .C (x2), .Y (n5994) );
  NOR2x1_ASAP7_75t_R   g5987( .A (n5994), .B (n1646), .Y (n5995) );
  AND3x1_ASAP7_75t_R   g5988( .A (n15), .B (x3), .C (x5), .Y (n5996) );
  NAND2x1_ASAP7_75t_R  g5989( .A (x4), .B (n5996), .Y (n5997) );
  INVx1_ASAP7_75t_R    g5990( .A (n5997), .Y (n5998) );
  AO21x1_ASAP7_75t_R   g5991( .A1 (n5993), .A2 (n5995), .B (n5998), .Y (y2834) );
  INVx1_ASAP7_75t_R    g5992( .A (n148), .Y (n6000) );
  AO21x1_ASAP7_75t_R   g5993( .A1 (n1564), .A2 (n63), .B (n6000), .Y (n6001) );
  OA21x2_ASAP7_75t_R   g5994( .A1 (n148), .A2 (n1590), .B (n6001), .Y (y2835) );
  AO21x1_ASAP7_75t_R   g5995( .A1 (y2079), .A2 (x4), .B (n300), .Y (y2836) );
  NAND2x1_ASAP7_75t_R  g5996( .A (x4), .B (n3645), .Y (n6004) );
  AO32x1_ASAP7_75t_R   g5997( .A1 (n17), .A2 (n556), .A3 (x0), .B1 (y2079), .B2 (n6004), .Y (y2837) );
  AND2x2_ASAP7_75t_R   g5998( .A (n1175), .B (y2079), .Y (y2838) );
  OR3x1_ASAP7_75t_R    g5999( .A (n3628), .B (n3490), .C (n1269), .Y (y2839) );
  AO21x1_ASAP7_75t_R   g6000( .A1 (n4057), .A2 (x3), .B (n4217), .Y (y2840) );
  OR3x1_ASAP7_75t_R    g6001( .A (n3399), .B (n306), .C (n354), .Y (y2841) );
  INVx1_ASAP7_75t_R    g6002( .A (n3445), .Y (n6010) );
  AO21x1_ASAP7_75t_R   g6003( .A1 (n316), .A2 (n15), .B (n3207), .Y (n6011) );
  OA21x2_ASAP7_75t_R   g6004( .A1 (n3963), .A2 (n6010), .B (n6011), .Y (y2842) );
  AO21x1_ASAP7_75t_R   g6005( .A1 (n17), .A2 (n4028), .B (n332), .Y (y2843) );
  INVx1_ASAP7_75t_R    g6006( .A (n3629), .Y (n6014) );
  AO32x1_ASAP7_75t_R   g6007( .A1 (n1265), .A2 (n293), .A3 (n3567), .B1 (n97), .B2 (n6014), .Y (y2844) );
  AO21x1_ASAP7_75t_R   g6008( .A1 (n3905), .A2 (n3278), .B (n5427), .Y (y2845) );
  OA21x2_ASAP7_75t_R   g6009( .A1 (n1775), .A2 (n1150), .B (n299), .Y (y2846) );
  AND3x1_ASAP7_75t_R   g6010( .A (n3380), .B (n219), .C (n455), .Y (y2847) );
  OR3x1_ASAP7_75t_R    g6011( .A (n337), .B (n12), .C (x5), .Y (n6019) );
  NAND2x1_ASAP7_75t_R  g6012( .A (n6019), .B (n3256), .Y (y2848) );
  INVx1_ASAP7_75t_R    g6013( .A (n3642), .Y (y2849) );
  AO21x1_ASAP7_75t_R   g6014( .A1 (n22), .A2 (n77), .B (n3963), .Y (y2887) );
  OA21x2_ASAP7_75t_R   g6015( .A1 (n3859), .A2 (n3282), .B (y2887), .Y (y2850) );
  OA21x2_ASAP7_75t_R   g6016( .A1 (n3568), .A2 (n3001), .B (n5688), .Y (y2851) );
  NOR2x1_ASAP7_75t_R   g6017( .A (n22), .B (n5543), .Y (n6025) );
  AO21x1_ASAP7_75t_R   g6018( .A1 (n3823), .A2 (n5370), .B (n6025), .Y (y2853) );
  NAND2x1_ASAP7_75t_R  g6019( .A (n1528), .B (n1527), .Y (y2854) );
  OA21x2_ASAP7_75t_R   g6020( .A1 (n492), .A2 (n994), .B (n1167), .Y (y2855) );
  AO21x1_ASAP7_75t_R   g6021( .A1 (n218), .A2 (n29), .B (n3963), .Y (y2856) );
  AO32x1_ASAP7_75t_R   g6022( .A1 (n22), .A2 (n97), .A3 (n316), .B1 (x4), .B2 (n5654), .Y (y2857) );
  OA22x2_ASAP7_75t_R   g6023( .A1 (n492), .A2 (n994), .B1 (n1775), .B2 (n970), .Y (y2858) );
  OR3x1_ASAP7_75t_R    g6024( .A (n186), .B (y863), .C (n856), .Y (y2859) );
  AO21x1_ASAP7_75t_R   g6025( .A1 (n316), .A2 (n319), .B (x2), .Y (n6033) );
  OA21x2_ASAP7_75t_R   g6026( .A1 (n3960), .A2 (n3025), .B (n6033), .Y (y2860) );
  NOR2x1_ASAP7_75t_R   g6027( .A (n352), .B (n436), .Y (n6035) );
  INVx1_ASAP7_75t_R    g6028( .A (n6035), .Y (n6036) );
  AND2x2_ASAP7_75t_R   g6029( .A (n6036), .B (n4357), .Y (y2861) );
  AND2x2_ASAP7_75t_R   g6030( .A (n4667), .B (y2079), .Y (y2862) );
  OA21x2_ASAP7_75t_R   g6031( .A1 (n3298), .A2 (n5108), .B (n3705), .Y (y2863) );
  AND3x1_ASAP7_75t_R   g6032( .A (n765), .B (n466), .C (n2008), .Y (n6040) );
  INVx1_ASAP7_75t_R    g6033( .A (n6040), .Y (n6041) );
  AND3x1_ASAP7_75t_R   g6034( .A (n6041), .B (n4083), .C (n556), .Y (y2864) );
  NOR2x1_ASAP7_75t_R   g6035( .A (n17), .B (n756), .Y (n6043) );
  AO21x1_ASAP7_75t_R   g6036( .A1 (x4), .A2 (n6043), .B (n4077), .Y (y2865) );
  AO21x1_ASAP7_75t_R   g6037( .A1 (n17), .A2 (x2), .B (y2079), .Y (n6045) );
  AO32x1_ASAP7_75t_R   g6038( .A1 (x3), .A2 (n3028), .A3 (x5), .B1 (n6045), .B2 (n360), .Y (y2866) );
  AND2x2_ASAP7_75t_R   g6039( .A (n2490), .B (n64), .Y (y2867) );
  NAND2x1_ASAP7_75t_R  g6040( .A (x2), .B (y2022), .Y (n6048) );
  INVx1_ASAP7_75t_R    g6041( .A (n6048), .Y (y2868) );
  AO21x1_ASAP7_75t_R   g6042( .A1 (n576), .A2 (n17), .B (n3234), .Y (y2869) );
  AO21x1_ASAP7_75t_R   g6043( .A1 (n1262), .A2 (n765), .B (n143), .Y (y2870) );
  OAI21x1_ASAP7_75t_R  g6044( .A1 (n3316), .A2 (n2997), .B (n28), .Y (y2871) );
  AND3x1_ASAP7_75t_R   g6045( .A (y2196), .B (n63), .C (n64), .Y (y2873) );
  AND2x2_ASAP7_75t_R   g6046( .A (y2305), .B (n453), .Y (y2874) );
  AND2x2_ASAP7_75t_R   g6047( .A (n4353), .B (n3119), .Y (y2875) );
  AO21x1_ASAP7_75t_R   g6048( .A1 (n5385), .A2 (x3), .B (n638), .Y (y2876) );
  AND2x2_ASAP7_75t_R   g6049( .A (n963), .B (n1077), .Y (y2877) );
  AND2x2_ASAP7_75t_R   g6050( .A (n3380), .B (n1272), .Y (y2879) );
  AND2x2_ASAP7_75t_R   g6051( .A (y1742), .B (x0), .Y (y2880) );
  INVx1_ASAP7_75t_R    g6052( .A (n724), .Y (n6060) );
  AO21x1_ASAP7_75t_R   g6053( .A1 (n3646), .A2 (x4), .B (n6060), .Y (n6061) );
  NOR2x1_ASAP7_75t_R   g6054( .A (n481), .B (n6061), .Y (y2881) );
  AND2x2_ASAP7_75t_R   g6055( .A (n3459), .B (n4341), .Y (y2883) );
  INVx1_ASAP7_75t_R    g6056( .A (n1253), .Y (n6064) );
  AND3x1_ASAP7_75t_R   g6057( .A (n6064), .B (n1295), .C (x2), .Y (n6065) );
  OA21x2_ASAP7_75t_R   g6058( .A1 (n2889), .A2 (n1253), .B (n15), .Y (n6066) );
  AO21x1_ASAP7_75t_R   g6059( .A1 (n16), .A2 (x3), .B (n12), .Y (n6067) );
  INVx1_ASAP7_75t_R    g6060( .A (n6067), .Y (n6068) );
  OR3x1_ASAP7_75t_R    g6061( .A (n6065), .B (n6066), .C (n6068), .Y (y2884) );
  AND2x2_ASAP7_75t_R   g6062( .A (n1863), .B (y1845), .Y (y2885) );
  OA21x2_ASAP7_75t_R   g6063( .A1 (n1223), .A2 (n4166), .B (y3293), .Y (y2886) );
  OA21x2_ASAP7_75t_R   g6064( .A1 (n3182), .A2 (n3918), .B (n5830), .Y (y2888) );
  AO21x1_ASAP7_75t_R   g6065( .A1 (y9), .A2 (n310), .B (n527), .Y (n6073) );
  OA21x2_ASAP7_75t_R   g6066( .A1 (x5), .A2 (n6073), .B (y2737), .Y (y2889) );
  AO21x1_ASAP7_75t_R   g6067( .A1 (n3866), .A2 (n3025), .B (n3819), .Y (y2890) );
  NAND2x1_ASAP7_75t_R  g6068( .A (n3083), .B (n5465), .Y (y2891) );
  AND2x2_ASAP7_75t_R   g6069( .A (n5435), .B (n5081), .Y (y2892) );
  AO21x1_ASAP7_75t_R   g6070( .A1 (n1540), .A2 (n228), .B (n2865), .Y (y2893) );
  AND3x1_ASAP7_75t_R   g6071( .A (y2196), .B (n360), .C (n290), .Y (n6079) );
  INVx1_ASAP7_75t_R    g6072( .A (n6079), .Y (n6080) );
  AND2x2_ASAP7_75t_R   g6073( .A (n6080), .B (y3198), .Y (y2894) );
  OR3x1_ASAP7_75t_R    g6074( .A (n4575), .B (n3447), .C (n4576), .Y (y2895) );
  OA211x2_ASAP7_75t_R  g6075( .A1 (n4916), .A2 (n4621), .B (n5109), .C (n556), .Y (y2896) );
  XNOR2x2_ASAP7_75t_R  g6076( .A (n1903), .B (n3093), .Y (y2897) );
  AO21x1_ASAP7_75t_R   g6077( .A1 (n173), .A2 (x5), .B (n3732), .Y (n6085) );
  NAND2x1_ASAP7_75t_R  g6078( .A (n1738), .B (n6085), .Y (y2898) );
  AO21x1_ASAP7_75t_R   g6079( .A1 (x4), .A2 (n12), .B (n369), .Y (n6087) );
  OA21x2_ASAP7_75t_R   g6080( .A1 (n29), .A2 (n5111), .B (n6087), .Y (y2899) );
  OA21x2_ASAP7_75t_R   g6081( .A1 (n4584), .A2 (y1300), .B (n1334), .Y (y2901) );
  AND3x1_ASAP7_75t_R   g6082( .A (n4109), .B (n4151), .C (n556), .Y (y2902) );
  OR3x1_ASAP7_75t_R    g6083( .A (n3112), .B (n22), .C (n3192), .Y (n6091) );
  AND2x2_ASAP7_75t_R   g6084( .A (n6091), .B (n5964), .Y (y2903) );
  NOR2x1_ASAP7_75t_R   g6085( .A (x5), .B (n3989), .Y (y2905) );
  AND3x1_ASAP7_75t_R   g6086( .A (n3797), .B (n3139), .C (n556), .Y (y2906) );
  AND2x2_ASAP7_75t_R   g6087( .A (y1693), .B (x0), .Y (y2907) );
  AND3x1_ASAP7_75t_R   g6088( .A (n3705), .B (n4151), .C (n556), .Y (y2908) );
  OR3x1_ASAP7_75t_R    g6089( .A (n4625), .B (y2022), .C (x2), .Y (n6097) );
  AND3x1_ASAP7_75t_R   g6090( .A (n6097), .B (n2307), .C (y3852), .Y (y2909) );
  AO21x1_ASAP7_75t_R   g6091( .A1 (n3023), .A2 (n3776), .B (n2964), .Y (y2910) );
  AND2x2_ASAP7_75t_R   g6092( .A (n4588), .B (n3919), .Y (y2911) );
  OR3x1_ASAP7_75t_R    g6093( .A (n5077), .B (n3634), .C (n3189), .Y (y2912) );
  AO21x1_ASAP7_75t_R   g6094( .A1 (n4804), .A2 (n77), .B (y2079), .Y (y2913) );
  INVx1_ASAP7_75t_R    g6095( .A (n4094), .Y (n6103) );
  OA21x2_ASAP7_75t_R   g6096( .A1 (n337), .A2 (n4022), .B (n6103), .Y (y2914) );
  NOR2x1_ASAP7_75t_R   g6097( .A (n2441), .B (n1527), .Y (n6105) );
  OA21x2_ASAP7_75t_R   g6098( .A1 (n6105), .A2 (x3), .B (n2552), .Y (y2915) );
  AO21x1_ASAP7_75t_R   g6099( .A1 (y2079), .A2 (n22), .B (n211), .Y (n6107) );
  INVx1_ASAP7_75t_R    g6100( .A (n6107), .Y (n6108) );
  INVx1_ASAP7_75t_R    g6101( .A (n3430), .Y (n6109) );
  AO21x1_ASAP7_75t_R   g6102( .A1 (n4633), .A2 (n6108), .B (n6109), .Y (y2917) );
  OR3x1_ASAP7_75t_R    g6103( .A (n29), .B (n2718), .C (n1775), .Y (y3269) );
  AO21x1_ASAP7_75t_R   g6104( .A1 (n28), .A2 (n614), .B (x3), .Y (n6112) );
  AND2x2_ASAP7_75t_R   g6105( .A (y3269), .B (n6112), .Y (y2918) );
  NAND2x1_ASAP7_75t_R  g6106( .A (n3040), .B (n285), .Y (y2919) );
  NOR2x1_ASAP7_75t_R   g6107( .A (x5), .B (n4439), .Y (n6115) );
  AO21x1_ASAP7_75t_R   g6108( .A1 (x5), .A2 (n4518), .B (n6115), .Y (n6116) );
  XOR2x2_ASAP7_75t_R   g6109( .A (n6116), .B (n17), .Y (y2920) );
  AO21x1_ASAP7_75t_R   g6110( .A1 (n144), .A2 (x2), .B (n1911), .Y (n6118) );
  AO21x1_ASAP7_75t_R   g6111( .A1 (n2116), .A2 (n2117), .B (n17), .Y (n6119) );
  OA21x2_ASAP7_75t_R   g6112( .A1 (n1295), .A2 (n6118), .B (n6119), .Y (y2921) );
  AO32x1_ASAP7_75t_R   g6113( .A1 (n17), .A2 (n5085), .A3 (n4056), .B1 (x3), .B2 (n4057), .Y (y2922) );
  NAND2x1_ASAP7_75t_R  g6114( .A (n137), .B (n28), .Y (n6122) );
  NAND2x1_ASAP7_75t_R  g6115( .A (n72), .B (n388), .Y (n6123) );
  XOR2x2_ASAP7_75t_R   g6116( .A (n6122), .B (n6123), .Y (y2923) );
  AO21x1_ASAP7_75t_R   g6117( .A1 (n90), .A2 (n219), .B (x4), .Y (n6125) );
  INVx1_ASAP7_75t_R    g6118( .A (n6125), .Y (n6126) );
  OR3x1_ASAP7_75t_R    g6119( .A (n6126), .B (n911), .C (n529), .Y (y2924) );
  INVx1_ASAP7_75t_R    g6120( .A (n3588), .Y (n6128) );
  OA21x2_ASAP7_75t_R   g6121( .A1 (n4373), .A2 (n6128), .B (y3397), .Y (y2925) );
  AO21x1_ASAP7_75t_R   g6122( .A1 (n22), .A2 (n3004), .B (n4554), .Y (y2926) );
  AO32x1_ASAP7_75t_R   g6123( .A1 (y2079), .A2 (n299), .A3 (n310), .B1 (x5), .B2 (n3267), .Y (n6131) );
  NAND2x1_ASAP7_75t_R  g6124( .A (n4635), .B (n6131), .Y (y2927) );
  OR3x1_ASAP7_75t_R    g6125( .A (n503), .B (n563), .C (n537), .Y (y2928) );
  AND3x1_ASAP7_75t_R   g6126( .A (n700), .B (n740), .C (n776), .Y (n6134) );
  OA21x2_ASAP7_75t_R   g6127( .A1 (x0), .A2 (n6134), .B (n1331), .Y (y2929) );
  AO32x1_ASAP7_75t_R   g6128( .A1 (y2079), .A2 (n401), .A3 (n72), .B1 (n3909), .B2 (n22), .Y (y2930) );
  NAND2x1_ASAP7_75t_R  g6129( .A (x2), .B (n349), .Y (n6137) );
  INVx1_ASAP7_75t_R    g6130( .A (n6137), .Y (n6138) );
  INVx1_ASAP7_75t_R    g6131( .A (n2979), .Y (n6139) );
  OR3x1_ASAP7_75t_R    g6132( .A (n6138), .B (n6139), .C (n347), .Y (y2931) );
  NAND2x1_ASAP7_75t_R  g6133( .A (n17), .B (n439), .Y (n6141) );
  OA21x2_ASAP7_75t_R   g6134( .A1 (n3116), .A2 (y2079), .B (n6141), .Y (y2932) );
  OA22x2_ASAP7_75t_R   g6135( .A1 (n3819), .A2 (n3618), .B1 (n1646), .B2 (n3181), .Y (y2933) );
  AND2x2_ASAP7_75t_R   g6136( .A (n3455), .B (n1272), .Y (y2934) );
  AO21x1_ASAP7_75t_R   g6137( .A1 (n5227), .A2 (n3284), .B (n5214), .Y (y2935) );
  AND2x2_ASAP7_75t_R   g6138( .A (y1227), .B (n4504), .Y (y2936) );
  AO21x1_ASAP7_75t_R   g6139( .A1 (y2079), .A2 (n3377), .B (n4230), .Y (y2937) );
  AO21x1_ASAP7_75t_R   g6140( .A1 (x3), .A2 (n1269), .B (n4964), .Y (y2938) );
  OA21x2_ASAP7_75t_R   g6141( .A1 (n403), .A2 (n4528), .B (y3397), .Y (y2939) );
  AO21x1_ASAP7_75t_R   g6142( .A1 (n17), .A2 (n3000), .B (n164), .Y (n6150) );
  INVx1_ASAP7_75t_R    g6143( .A (n6150), .Y (n6151) );
  AO21x1_ASAP7_75t_R   g6144( .A1 (n6151), .A2 (y2079), .B (n3525), .Y (y2940) );
  AND2x2_ASAP7_75t_R   g6145( .A (n5132), .B (n3256), .Y (y2941) );
  AND2x2_ASAP7_75t_R   g6146( .A (n2699), .B (n1772), .Y (y2942) );
  OA211x2_ASAP7_75t_R  g6147( .A1 (n369), .A2 (n2999), .B (n4536), .C (n1265), .Y (y2943) );
  AND3x1_ASAP7_75t_R   g6148( .A (n2322), .B (n2116), .C (n244), .Y (y2944) );
  INVx1_ASAP7_75t_R    g6149( .A (n632), .Y (n6157) );
  AO21x1_ASAP7_75t_R   g6150( .A1 (n5438), .A2 (x3), .B (n6157), .Y (n6158) );
  NAND2x1_ASAP7_75t_R  g6151( .A (n292), .B (n3457), .Y (n6159) );
  AND2x2_ASAP7_75t_R   g6152( .A (n6159), .B (x2), .Y (n6160) );
  AO21x1_ASAP7_75t_R   g6153( .A1 (n15), .A2 (n6158), .B (n6160), .Y (y2945) );
  OR3x1_ASAP7_75t_R    g6154( .A (n403), .B (y2079), .C (x2), .Y (n6162) );
  INVx1_ASAP7_75t_R    g6155( .A (n6162), .Y (n6163) );
  OR3x1_ASAP7_75t_R    g6156( .A (n6163), .B (n3611), .C (n337), .Y (y2946) );
  AND3x1_ASAP7_75t_R   g6157( .A (n4171), .B (n4341), .C (n72), .Y (y2947) );
  AND2x2_ASAP7_75t_R   g6158( .A (n5768), .B (n762), .Y (y2948) );
  AO21x1_ASAP7_75t_R   g6159( .A1 (n4336), .A2 (n3415), .B (n4349), .Y (y2949) );
  AND3x1_ASAP7_75t_R   g6160( .A (n4647), .B (n4089), .C (n4638), .Y (y2950) );
  AND2x2_ASAP7_75t_R   g6161( .A (n4504), .B (y1474), .Y (y2951) );
  AO21x1_ASAP7_75t_R   g6162( .A1 (n2790), .A2 (n1698), .B (n81), .Y (n6170) );
  AND2x2_ASAP7_75t_R   g6163( .A (n6170), .B (n219), .Y (y2952) );
  AND3x1_ASAP7_75t_R   g6164( .A (n337), .B (y2079), .C (x0), .Y (y3262) );
  INVx1_ASAP7_75t_R    g6165( .A (y3262), .Y (n6173) );
  INVx1_ASAP7_75t_R    g6166( .A (n4478), .Y (n6174) );
  AND3x1_ASAP7_75t_R   g6167( .A (n6173), .B (y1702), .C (n6174), .Y (y2953) );
  INVx1_ASAP7_75t_R    g6168( .A (n4586), .Y (n6176) );
  AND3x1_ASAP7_75t_R   g6169( .A (n6176), .B (n366), .C (x2), .Y (n6177) );
  AO21x1_ASAP7_75t_R   g6170( .A1 (n650), .A2 (n3144), .B (n6177), .Y (y2954) );
  OA21x2_ASAP7_75t_R   g6171( .A1 (n4313), .A2 (n700), .B (n3712), .Y (y2955) );
  AND3x1_ASAP7_75t_R   g6172( .A (n4111), .B (n5435), .C (y1281), .Y (y2956) );
  AO21x1_ASAP7_75t_R   g6173( .A1 (n22), .A2 (n3828), .B (n3611), .Y (y2957) );
  OR3x1_ASAP7_75t_R    g6174( .A (n628), .B (n3568), .C (n3263), .Y (y2958) );
  AND3x1_ASAP7_75t_R   g6175( .A (n4317), .B (n3023), .C (n5507), .Y (y2959) );
  AND2x2_ASAP7_75t_R   g6176( .A (y2727), .B (n3648), .Y (y2960) );
  AO21x1_ASAP7_75t_R   g6177( .A1 (n72), .A2 (n137), .B (y2079), .Y (n6185) );
  INVx1_ASAP7_75t_R    g6178( .A (n6185), .Y (n6186) );
  INVx1_ASAP7_75t_R    g6179( .A (n5128), .Y (n6187) );
  OA21x2_ASAP7_75t_R   g6180( .A1 (n6186), .A2 (n6187), .B (n556), .Y (y2961) );
  OR3x1_ASAP7_75t_R    g6181( .A (n3899), .B (n3132), .C (n81), .Y (y2962) );
  NAND2x1_ASAP7_75t_R  g6182( .A (n28), .B (n290), .Y (n6190) );
  AO21x1_ASAP7_75t_R   g6183( .A1 (n6190), .A2 (n15), .B (n5809), .Y (y2963) );
  AO21x1_ASAP7_75t_R   g6184( .A1 (n4588), .A2 (n22), .B (n5633), .Y (n6192) );
  AND2x2_ASAP7_75t_R   g6185( .A (n6192), .B (n5939), .Y (y2964) );
  AO21x1_ASAP7_75t_R   g6186( .A1 (n4089), .A2 (n2998), .B (n81), .Y (y2965) );
  AO21x1_ASAP7_75t_R   g6187( .A1 (n3629), .A2 (n3630), .B (n3628), .Y (y2966) );
  AO21x1_ASAP7_75t_R   g6188( .A1 (n3457), .A2 (n292), .B (x2), .Y (n6196) );
  OA21x2_ASAP7_75t_R   g6189( .A1 (y1786), .A2 (n15), .B (n6196), .Y (y2967) );
  AO21x1_ASAP7_75t_R   g6190( .A1 (n22), .A2 (n17), .B (n756), .Y (n6198) );
  INVx1_ASAP7_75t_R    g6191( .A (n4514), .Y (n6199) );
  OAI21x1_ASAP7_75t_R  g6192( .A1 (n3310), .A2 (n6198), .B (n6199), .Y (y2968) );
  AO21x1_ASAP7_75t_R   g6193( .A1 (n1082), .A2 (x0), .B (n1924), .Y (y2969) );
  NAND2x1_ASAP7_75t_R  g6194( .A (n4233), .B (n382), .Y (n6202) );
  AOI21x1_ASAP7_75t_R  g6195( .A1 (n740), .A2 (n6202), .B (n5994), .Y (y2970) );
  AO21x1_ASAP7_75t_R   g6196( .A1 (n6199), .A2 (n5243), .B (n325), .Y (n6204) );
  NAND2x1_ASAP7_75t_R  g6197( .A (n740), .B (n6204), .Y (y2971) );
  AND2x2_ASAP7_75t_R   g6198( .A (n2980), .B (x5), .Y (n6206) );
  OAI21x1_ASAP7_75t_R  g6199( .A1 (n6206), .A2 (n3608), .B (n348), .Y (y2972) );
  INVx1_ASAP7_75t_R    g6200( .A (n214), .Y (y2973) );
  OA21x2_ASAP7_75t_R   g6201( .A1 (n3580), .A2 (n4269), .B (y1903), .Y (y2974) );
  AND2x2_ASAP7_75t_R   g6202( .A (y1267), .B (n4638), .Y (y2975) );
  NAND2x1_ASAP7_75t_R  g6203( .A (n1186), .B (n697), .Y (y2976) );
  NAND2x1_ASAP7_75t_R  g6204( .A (x2), .B (n611), .Y (n6212) );
  AND2x2_ASAP7_75t_R   g6205( .A (n6212), .B (n2728), .Y (y2977) );
  OA33x2_ASAP7_75t_R   g6206( .A1 (n3027), .A2 (n17), .A3 (n5690), .B1 (y2079), .B2 (n3637), .B3 (n3568), .Y (y2978) );
  AO21x1_ASAP7_75t_R   g6207( .A1 (n700), .A2 (n707), .B (n2090), .Y (y2979) );
  AO21x1_ASAP7_75t_R   g6208( .A1 (n1510), .A2 (x0), .B (n53), .Y (y2980) );
  AO21x1_ASAP7_75t_R   g6209( .A1 (n4070), .A2 (n2971), .B (n3899), .Y (y2981) );
  INVx1_ASAP7_75t_R    g6210( .A (n3184), .Y (n6218) );
  OR3x1_ASAP7_75t_R    g6211( .A (n529), .B (n29), .C (n6218), .Y (y3387) );
  AO21x1_ASAP7_75t_R   g6212( .A1 (n388), .A2 (n28), .B (x2), .Y (n6220) );
  AND2x2_ASAP7_75t_R   g6213( .A (y3387), .B (n6220), .Y (y2982) );
  AND2x2_ASAP7_75t_R   g6214( .A (n2522), .B (n2532), .Y (y2983) );
  AO21x1_ASAP7_75t_R   g6215( .A1 (x4), .A2 (x5), .B (n211), .Y (n6223) );
  AND2x2_ASAP7_75t_R   g6216( .A (y1287), .B (n6223), .Y (y2984) );
  AND2x2_ASAP7_75t_R   g6217( .A (y1393), .B (n906), .Y (y2985) );
  AND2x2_ASAP7_75t_R   g6218( .A (n3395), .B (n463), .Y (y2986) );
  OA21x2_ASAP7_75t_R   g6219( .A1 (n396), .A2 (n211), .B (y1287), .Y (y2987) );
  INVx1_ASAP7_75t_R    g6220( .A (n5800), .Y (n6228) );
  NAND2x1_ASAP7_75t_R  g6221( .A (n17), .B (n5296), .Y (n6229) );
  INVx1_ASAP7_75t_R    g6222( .A (n6229), .Y (n6230) );
  OA21x2_ASAP7_75t_R   g6223( .A1 (n6228), .A2 (n6230), .B (n3011), .Y (y2988) );
  OA21x2_ASAP7_75t_R   g6224( .A1 (n389), .A2 (n4754), .B (n5484), .Y (y2989) );
  AND2x2_ASAP7_75t_R   g6225( .A (n97), .B (n740), .Y (n6233) );
  INVx1_ASAP7_75t_R    g6226( .A (n6233), .Y (n6234) );
  AND2x2_ASAP7_75t_R   g6227( .A (n97), .B (n360), .Y (n6235) );
  INVx1_ASAP7_75t_R    g6228( .A (n6235), .Y (n6236) );
  AO21x1_ASAP7_75t_R   g6229( .A1 (n97), .A2 (n740), .B (n291), .Y (n6237) );
  AO32x1_ASAP7_75t_R   g6230( .A1 (n290), .A2 (n6234), .A3 (n6235), .B1 (n6236), .B2 (n6237), .Y (y2990) );
  NAND2x1_ASAP7_75t_R  g6231( .A (n15), .B (n3565), .Y (n6239) );
  INVx1_ASAP7_75t_R    g6232( .A (n6239), .Y (n6240) );
  AO21x1_ASAP7_75t_R   g6233( .A1 (x5), .A2 (n4518), .B (n628), .Y (n6241) );
  AO21x1_ASAP7_75t_R   g6234( .A1 (n6240), .A2 (x4), .B (n6241), .Y (y2992) );
  OR3x1_ASAP7_75t_R    g6235( .A (n2202), .B (n1503), .C (n1269), .Y (y2993) );
  OA21x2_ASAP7_75t_R   g6236( .A1 (n15), .A2 (y1356), .B (n1912), .Y (y2994) );
  AO21x1_ASAP7_75t_R   g6237( .A1 (n1997), .A2 (x0), .B (y2466), .Y (n6245) );
  AND2x2_ASAP7_75t_R   g6238( .A (n6245), .B (n3119), .Y (y2995) );
  NAND2x1_ASAP7_75t_R  g6239( .A (n15), .B (y195), .Y (n6247) );
  AO32x1_ASAP7_75t_R   g6240( .A1 (y2079), .A2 (n6247), .A3 (n187), .B1 (x0), .B2 (n1643), .Y (y2996) );
  AO21x1_ASAP7_75t_R   g6241( .A1 (n1939), .A2 (n382), .B (x2), .Y (n6249) );
  OA21x2_ASAP7_75t_R   g6242( .A1 (y1445), .A2 (n15), .B (n6249), .Y (y2997) );
  AO21x1_ASAP7_75t_R   g6243( .A1 (x5), .A2 (n3263), .B (n4991), .Y (y2998) );
  AO21x1_ASAP7_75t_R   g6244( .A1 (n17), .A2 (x0), .B (x5), .Y (n6252) );
  INVx1_ASAP7_75t_R    g6245( .A (n6252), .Y (n6253) );
  OR3x1_ASAP7_75t_R    g6246( .A (n1158), .B (n291), .C (n6253), .Y (n6254) );
  AND2x2_ASAP7_75t_R   g6247( .A (n6254), .B (n3477), .Y (y2999) );
  OR3x1_ASAP7_75t_R    g6248( .A (n315), .B (x5), .C (x3), .Y (n6256) );
  OA21x2_ASAP7_75t_R   g6249( .A1 (n5633), .A2 (n3414), .B (n6256), .Y (y3000) );
  AND3x1_ASAP7_75t_R   g6250( .A (n388), .B (n28), .C (n15), .Y (n6258) );
  INVx1_ASAP7_75t_R    g6251( .A (n6258), .Y (n6259) );
  AND2x2_ASAP7_75t_R   g6252( .A (n3297), .B (x3), .Y (n6260) );
  AOI21x1_ASAP7_75t_R  g6253( .A1 (n17), .A2 (n6259), .B (n6260), .Y (y3002) );
  AO21x1_ASAP7_75t_R   g6254( .A1 (n1046), .A2 (n219), .B (n344), .Y (y3003) );
  OA21x2_ASAP7_75t_R   g6255( .A1 (n1054), .A2 (y1850), .B (n1023), .Y (y3004) );
  INVx1_ASAP7_75t_R    g6256( .A (n3443), .Y (n6264) );
  AO21x1_ASAP7_75t_R   g6257( .A1 (n22), .A2 (x5), .B (n3443), .Y (n6265) );
  AO32x1_ASAP7_75t_R   g6258( .A1 (n28), .A2 (n6264), .A3 (x2), .B1 (n15), .B2 (n6265), .Y (n6266) );
  NOR2x1_ASAP7_75t_R   g6259( .A (n218), .B (n6266), .Y (y3005) );
  XNOR2x2_ASAP7_75t_R  g6260( .A (n2992), .B (n5633), .Y (y3006) );
  INVx1_ASAP7_75t_R    g6261( .A (n2254), .Y (n6269) );
  OR3x1_ASAP7_75t_R    g6262( .A (n6269), .B (n619), .C (n276), .Y (y3007) );
  AO21x1_ASAP7_75t_R   g6263( .A1 (n316), .A2 (n319), .B (x4), .Y (n6271) );
  AO21x1_ASAP7_75t_R   g6264( .A1 (x3), .A2 (y2079), .B (n3028), .Y (n6272) );
  AND3x1_ASAP7_75t_R   g6265( .A (n6271), .B (n6272), .C (n72), .Y (y3008) );
  NAND2x1_ASAP7_75t_R  g6266( .A (n22), .B (n3588), .Y (n6274) );
  AO21x1_ASAP7_75t_R   g6267( .A1 (n15), .A2 (n17), .B (n3611), .Y (n6275) );
  OAI21x1_ASAP7_75t_R  g6268( .A1 (n6274), .A2 (n6275), .B (n3613), .Y (y3009) );
  AO21x1_ASAP7_75t_R   g6269( .A1 (n3612), .A2 (n3588), .B (x4), .Y (n6277) );
  OR3x1_ASAP7_75t_R    g6270( .A (n3611), .B (n22), .C (n45), .Y (n6278) );
  AND2x2_ASAP7_75t_R   g6271( .A (n6277), .B (n6278), .Y (y3010) );
  NOR2x1_ASAP7_75t_R   g6272( .A (n918), .B (n3461), .Y (y3011) );
  AO21x1_ASAP7_75t_R   g6273( .A1 (n3298), .A2 (x3), .B (n3263), .Y (y3012) );
  AO21x1_ASAP7_75t_R   g6274( .A1 (n22), .A2 (n312), .B (n563), .Y (n6282) );
  AO21x1_ASAP7_75t_R   g6275( .A1 (n6282), .A2 (n497), .B (n537), .Y (y3013) );
  AO32x1_ASAP7_75t_R   g6276( .A1 (y2079), .A2 (n3448), .A3 (n4142), .B1 (n4495), .B2 (n4494), .Y (y3014) );
  AND2x2_ASAP7_75t_R   g6277( .A (n3457), .B (x2), .Y (n6285) );
  AO21x1_ASAP7_75t_R   g6278( .A1 (n6285), .A2 (n556), .B (n3263), .Y (y3015) );
  INVx1_ASAP7_75t_R    g6279( .A (n3278), .Y (n6287) );
  AO32x1_ASAP7_75t_R   g6280( .A1 (n1158), .A2 (n97), .A3 (n6287), .B1 (n3905), .B2 (n3278), .Y (y3016) );
  NAND2x1_ASAP7_75t_R  g6281( .A (n5109), .B (n3613), .Y (y3017) );
  AND2x2_ASAP7_75t_R   g6282( .A (n3681), .B (y3293), .Y (y3018) );
  AO21x1_ASAP7_75t_R   g6283( .A1 (n22), .A2 (x5), .B (x2), .Y (n6291) );
  INVx1_ASAP7_75t_R    g6284( .A (n6291), .Y (n6292) );
  INVx1_ASAP7_75t_R    g6285( .A (n5801), .Y (n6293) );
  OA22x2_ASAP7_75t_R   g6286( .A1 (n5801), .A2 (n6292), .B1 (n6293), .B2 (n5539), .Y (y3019) );
  NAND2x1_ASAP7_75t_R  g6287( .A (n12), .B (n1403), .Y (n6295) );
  AND2x2_ASAP7_75t_R   g6288( .A (n2639), .B (n6295), .Y (y3020) );
  AO21x1_ASAP7_75t_R   g6289( .A1 (y2740), .A2 (x0), .B (n2600), .Y (y3021) );
  AO32x1_ASAP7_75t_R   g6290( .A1 (x4), .A2 (n5176), .A3 (n6234), .B1 (n5177), .B2 (n4621), .Y (y3022) );
  OA21x2_ASAP7_75t_R   g6291( .A1 (n4631), .A2 (n418), .B (n3170), .Y (y3023) );
  OA21x2_ASAP7_75t_R   g6292( .A1 (n218), .A2 (n3446), .B (n3987), .Y (y3024) );
  AO21x1_ASAP7_75t_R   g6293( .A1 (x4), .A2 (n3294), .B (n1269), .Y (n6301) );
  AO32x1_ASAP7_75t_R   g6294( .A1 (n97), .A2 (n740), .A3 (n1158), .B1 (n4109), .B2 (n6301), .Y (y3025) );
  AO21x1_ASAP7_75t_R   g6295( .A1 (n3474), .A2 (x0), .B (n5271), .Y (y3026) );
  NAND2x1_ASAP7_75t_R  g6296( .A (n28), .B (n125), .Y (n6304) );
  OA21x2_ASAP7_75t_R   g6297( .A1 (n6304), .A2 (n3443), .B (n4835), .Y (y3027) );
  INVx1_ASAP7_75t_R    g6298( .A (n4708), .Y (n6306) );
  AO21x1_ASAP7_75t_R   g6299( .A1 (n3568), .A2 (x3), .B (y2079), .Y (n6307) );
  AO21x1_ASAP7_75t_R   g6300( .A1 (n6306), .A2 (n15), .B (n6307), .Y (n6308) );
  AND2x2_ASAP7_75t_R   g6301( .A (n6308), .B (n3706), .Y (y3028) );
  OR3x1_ASAP7_75t_R    g6302( .A (n1646), .B (n1269), .C (n22), .Y (n6310) );
  AND3x1_ASAP7_75t_R   g6303( .A (n6310), .B (n72), .C (n401), .Y (y3029) );
  AO21x1_ASAP7_75t_R   g6304( .A1 (n369), .A2 (n1163), .B (n5111), .Y (y3030) );
  AO21x1_ASAP7_75t_R   g6305( .A1 (y9), .A2 (n556), .B (n143), .Y (n6313) );
  AO21x1_ASAP7_75t_R   g6306( .A1 (n3203), .A2 (n16), .B (n6313), .Y (y3031) );
  AND2x2_ASAP7_75t_R   g6307( .A (n2256), .B (n271), .Y (n6315) );
  AO21x1_ASAP7_75t_R   g6308( .A1 (x2), .A2 (n1668), .B (n6315), .Y (y3032) );
  AO21x1_ASAP7_75t_R   g6309( .A1 (n52), .A2 (n363), .B (y2259), .Y (y3033) );
  OA211x2_ASAP7_75t_R  g6310( .A1 (n3123), .A2 (x3), .B (n6310), .C (n72), .Y (y3034) );
  AND2x2_ASAP7_75t_R   g6311( .A (n6103), .B (n4022), .Y (y3035) );
  AO21x1_ASAP7_75t_R   g6312( .A1 (n97), .A2 (y752), .B (n2126), .Y (y3036) );
  AND3x1_ASAP7_75t_R   g6313( .A (n97), .B (n64), .C (n219), .Y (y3037) );
  OR3x1_ASAP7_75t_R    g6314( .A (n17), .B (y2079), .C (x2), .Y (n6322) );
  AO21x1_ASAP7_75t_R   g6315( .A1 (n5085), .A2 (n6322), .B (n1269), .Y (n6323) );
  AND2x2_ASAP7_75t_R   g6316( .A (n6323), .B (n401), .Y (y3038) );
  AND2x2_ASAP7_75t_R   g6317( .A (n3464), .B (n1265), .Y (y3039) );
  AO21x1_ASAP7_75t_R   g6318( .A1 (n1062), .A2 (x5), .B (n856), .Y (n6326) );
  AOI22x1_ASAP7_75t_R  g6319( .A1 (n3124), .A2 (n1838), .B1 (n6326), .B2 (x4), .Y (y3040) );
  OR3x1_ASAP7_75t_R    g6320( .A (n3296), .B (n5427), .C (n1269), .Y (y3041) );
  AND2x2_ASAP7_75t_R   g6321( .A (n770), .B (x0), .Y (n6329) );
  AO21x1_ASAP7_75t_R   g6322( .A1 (n750), .A2 (n752), .B (n6329), .Y (y3042) );
  INVx1_ASAP7_75t_R    g6323( .A (n3359), .Y (n6331) );
  OA21x2_ASAP7_75t_R   g6324( .A1 (n6331), .A2 (n638), .B (n388), .Y (n6332) );
  NOR2x1_ASAP7_75t_R   g6325( .A (n164), .B (n6332), .Y (y3043) );
  AO21x1_ASAP7_75t_R   g6326( .A1 (y2079), .A2 (x3), .B (n756), .Y (n6334) );
  AO21x1_ASAP7_75t_R   g6327( .A1 (n22), .A2 (n6334), .B (n4841), .Y (y3044) );
  AO21x1_ASAP7_75t_R   g6328( .A1 (n17), .A2 (x4), .B (n756), .Y (n6336) );
  NOR2x1_ASAP7_75t_R   g6329( .A (x5), .B (n4495), .Y (n6337) );
  AO21x1_ASAP7_75t_R   g6330( .A1 (n4495), .A2 (n6336), .B (n6337), .Y (y3045) );
  OR3x1_ASAP7_75t_R    g6331( .A (n3568), .B (n3443), .C (n45), .Y (y3046) );
  AND2x2_ASAP7_75t_R   g6332( .A (n2971), .B (n4638), .Y (n6340) );
  NOR2x1_ASAP7_75t_R   g6333( .A (n81), .B (n28), .Y (n6341) );
  AO21x1_ASAP7_75t_R   g6334( .A1 (n6340), .A2 (n3282), .B (n6341), .Y (y3048) );
  NAND2x1_ASAP7_75t_R  g6335( .A (n17), .B (n718), .Y (n6343) );
  AO21x1_ASAP7_75t_R   g6336( .A1 (n660), .A2 (y3852), .B (y2196), .Y (n6344) );
  OA21x2_ASAP7_75t_R   g6337( .A1 (n450), .A2 (n6343), .B (n6344), .Y (y3049) );
  AND3x1_ASAP7_75t_R   g6338( .A (n2882), .B (n152), .C (n1482), .Y (y3050) );
  NAND2x1_ASAP7_75t_R  g6339( .A (n43), .B (n740), .Y (y3939) );
  INVx1_ASAP7_75t_R    g6340( .A (y3939), .Y (n6348) );
  NOR2x1_ASAP7_75t_R   g6341( .A (n43), .B (n740), .Y (n6349) );
  OR3x1_ASAP7_75t_R    g6342( .A (n6348), .B (n6349), .C (n143), .Y (y3051) );
  NAND2x1_ASAP7_75t_R  g6343( .A (x3), .B (n4753), .Y (n6351) );
  AND2x2_ASAP7_75t_R   g6344( .A (n6103), .B (n6351), .Y (y3052) );
  AND2x2_ASAP7_75t_R   g6345( .A (y168), .B (n632), .Y (y3053) );
  OR3x1_ASAP7_75t_R    g6346( .A (n529), .B (n4576), .C (n3447), .Y (y3054) );
  OA22x2_ASAP7_75t_R   g6347( .A1 (n3123), .A2 (n2965), .B1 (n3278), .B2 (n22), .Y (y3055) );
  AND3x1_ASAP7_75t_R   g6348( .A (n3804), .B (n4070), .C (y2079), .Y (y3056) );
  AND2x2_ASAP7_75t_R   g6349( .A (n4341), .B (n72), .Y (n6357) );
  OA21x2_ASAP7_75t_R   g6350( .A1 (n3123), .A2 (x3), .B (n6357), .Y (y3057) );
  AO21x1_ASAP7_75t_R   g6351( .A1 (x3), .A2 (n537), .B (n337), .Y (n6359) );
  AND2x2_ASAP7_75t_R   g6352( .A (n6359), .B (y2079), .Y (n6360) );
  AO21x1_ASAP7_75t_R   g6353( .A1 (n2050), .A2 (x0), .B (n6360), .Y (y3058) );
  AND3x1_ASAP7_75t_R   g6354( .A (n3459), .B (n4341), .C (n401), .Y (y3059) );
  AND3x1_ASAP7_75t_R   g6355( .A (n3805), .B (n5910), .C (n3282), .Y (y3060) );
  AND2x2_ASAP7_75t_R   g6356( .A (y1903), .B (n4362), .Y (y3061) );
  AO21x1_ASAP7_75t_R   g6357( .A1 (n1572), .A2 (n360), .B (n2999), .Y (n6365) );
  AO21x1_ASAP7_75t_R   g6358( .A1 (y2079), .A2 (n6365), .B (n4878), .Y (y3062) );
  NOR2x1_ASAP7_75t_R   g6359( .A (y1281), .B (n3325), .Y (n6367) );
  AND2x2_ASAP7_75t_R   g6360( .A (y1281), .B (n3325), .Y (n6368) );
  OR3x1_ASAP7_75t_R    g6361( .A (n6367), .B (n6368), .C (y2466), .Y (y3063) );
  AND2x2_ASAP7_75t_R   g6362( .A (n3724), .B (y1871), .Y (y3064) );
  INVx1_ASAP7_75t_R    g6363( .A (n2998), .Y (n6371) );
  OR3x1_ASAP7_75t_R    g6364( .A (n6371), .B (y2079), .C (n3447), .Y (n6372) );
  OR3x1_ASAP7_75t_R    g6365( .A (n76), .B (n22), .C (x5), .Y (n6373) );
  AND3x1_ASAP7_75t_R   g6366( .A (n6372), .B (n6373), .C (n1572), .Y (y3065) );
  INVx1_ASAP7_75t_R    g6367( .A (n3832), .Y (n6375) );
  OA21x2_ASAP7_75t_R   g6368( .A1 (n4047), .A2 (n6375), .B (y3293), .Y (y3066) );
  AO21x1_ASAP7_75t_R   g6369( .A1 (n474), .A2 (n3191), .B (n529), .Y (y3067) );
  AND3x1_ASAP7_75t_R   g6370( .A (n3493), .B (n388), .C (n28), .Y (n6378) );
  AO21x1_ASAP7_75t_R   g6371( .A1 (y3758), .A2 (n3492), .B (n6378), .Y (n6379) );
  OR3x1_ASAP7_75t_R    g6372( .A (n6379), .B (n5665), .C (n347), .Y (y3068) );
  AND2x2_ASAP7_75t_R   g6373( .A (n5879), .B (n4904), .Y (y3069) );
  AO21x1_ASAP7_75t_R   g6374( .A1 (n718), .A2 (x3), .B (n3399), .Y (n6382) );
  AND2x2_ASAP7_75t_R   g6375( .A (n6382), .B (y3852), .Y (y3070) );
  AO21x1_ASAP7_75t_R   g6376( .A1 (n3023), .A2 (n3776), .B (n5858), .Y (y3071) );
  AND3x1_ASAP7_75t_R   g6377( .A (y2079), .B (n12), .C (x3), .Y (n6385) );
  AO21x1_ASAP7_75t_R   g6378( .A1 (x4), .A2 (n6385), .B (n5331), .Y (y3072) );
  AO21x1_ASAP7_75t_R   g6379( .A1 (n28), .A2 (n45), .B (n2989), .Y (n6387) );
  AO21x1_ASAP7_75t_R   g6380( .A1 (x4), .A2 (y2079), .B (n6387), .Y (y3073) );
  AND2x2_ASAP7_75t_R   g6381( .A (n4203), .B (y2648), .Y (y3075) );
  INVx1_ASAP7_75t_R    g6382( .A (n3083), .Y (n6390) );
  AO32x1_ASAP7_75t_R   g6383( .A1 (n22), .A2 (n3493), .A3 (n3083), .B1 (n6390), .B2 (n5465), .Y (y3076) );
  AND2x2_ASAP7_75t_R   g6384( .A (n5879), .B (n3000), .Y (y3077) );
  AO21x1_ASAP7_75t_R   g6385( .A1 (n1087), .A2 (n765), .B (n143), .Y (n6393) );
  AO21x1_ASAP7_75t_R   g6386( .A1 (n4028), .A2 (n352), .B (n6393), .Y (y3078) );
  OAI21x1_ASAP7_75t_R  g6387( .A1 (x5), .A2 (n1158), .B (n4465), .Y (y3079) );
  NOR2x1_ASAP7_75t_R   g6388( .A (n15), .B (n3118), .Y (n6396) );
  AO21x1_ASAP7_75t_R   g6389( .A1 (n396), .A2 (n164), .B (n6396), .Y (y3080) );
  INVx1_ASAP7_75t_R    g6390( .A (y2022), .Y (n6398) );
  AO21x1_ASAP7_75t_R   g6391( .A1 (n6398), .A2 (y9), .B (n1269), .Y (y3081) );
  NAND2x1_ASAP7_75t_R  g6392( .A (n3866), .B (n4465), .Y (y3082) );
  AO21x1_ASAP7_75t_R   g6393( .A1 (y2079), .A2 (x1), .B (n43), .Y (n6401) );
  NAND2x1_ASAP7_75t_R  g6394( .A (n2059), .B (n6401), .Y (y3083) );
  AO21x1_ASAP7_75t_R   g6395( .A1 (n15), .A2 (n17), .B (n518), .Y (n6403) );
  INVx1_ASAP7_75t_R    g6396( .A (n6403), .Y (n6404) );
  INVx1_ASAP7_75t_R    g6397( .A (n5701), .Y (n6405) );
  AO21x1_ASAP7_75t_R   g6398( .A1 (n3457), .A2 (n6404), .B (n6405), .Y (y3086) );
  INVx1_ASAP7_75t_R    g6399( .A (n2040), .Y (n6407) );
  AO21x1_ASAP7_75t_R   g6400( .A1 (y873), .A2 (x2), .B (n6407), .Y (y3087) );
  AND3x1_ASAP7_75t_R   g6401( .A (n583), .B (n369), .C (n290), .Y (y3088) );
  AND3x1_ASAP7_75t_R   g6402( .A (n5889), .B (n137), .C (n419), .Y (y3089) );
  OA211x2_ASAP7_75t_R  g6403( .A1 (n4526), .A2 (n5314), .B (n5484), .C (n72), .Y (y3090) );
  OA21x2_ASAP7_75t_R   g6404( .A1 (n529), .A2 (n442), .B (n219), .Y (y3091) );
  AO21x1_ASAP7_75t_R   g6405( .A1 (n295), .A2 (x2), .B (n164), .Y (n6413) );
  INVx1_ASAP7_75t_R    g6406( .A (n6413), .Y (y3092) );
  NOR2x1_ASAP7_75t_R   g6407( .A (n865), .B (n43), .Y (n6415) );
  AO21x1_ASAP7_75t_R   g6408( .A1 (x2), .A2 (n2565), .B (n6415), .Y (y3093) );
  AND3x1_ASAP7_75t_R   g6409( .A (n1272), .B (n1218), .C (n556), .Y (y3094) );
  AND3x1_ASAP7_75t_R   g6410( .A (y3293), .B (n391), .C (x2), .Y (n6418) );
  AO21x1_ASAP7_75t_R   g6411( .A1 (n419), .A2 (n45), .B (n6418), .Y (y3095) );
  AND2x2_ASAP7_75t_R   g6412( .A (n391), .B (x2), .Y (n6420) );
  AO21x1_ASAP7_75t_R   g6413( .A1 (n6420), .A2 (y3293), .B (n45), .Y (y3096) );
  INVx1_ASAP7_75t_R    g6414( .A (n1774), .Y (n6422) );
  OA21x2_ASAP7_75t_R   g6415( .A1 (n1064), .A2 (n6422), .B (y608), .Y (y3097) );
  AND2x2_ASAP7_75t_R   g6416( .A (y3198), .B (n299), .Y (y3098) );
  AO21x1_ASAP7_75t_R   g6417( .A1 (n22), .A2 (n1062), .B (n421), .Y (n6425) );
  AND3x1_ASAP7_75t_R   g6418( .A (n756), .B (n17), .C (n22), .Y (n6426) );
  INVx1_ASAP7_75t_R    g6419( .A (n6426), .Y (n6427) );
  AO21x1_ASAP7_75t_R   g6420( .A1 (n6425), .A2 (n6427), .B (n529), .Y (y3099) );
  OA21x2_ASAP7_75t_R   g6421( .A1 (n1458), .A2 (n826), .B (x5), .Y (n6429) );
  AOI21x1_ASAP7_75t_R  g6422( .A1 (n16), .A2 (n2060), .B (n6429), .Y (y3101) );
  OA21x2_ASAP7_75t_R   g6423( .A1 (n3027), .A2 (n4494), .B (n3302), .Y (y3102) );
  AND2x2_ASAP7_75t_R   g6424( .A (y1903), .B (n3326), .Y (y3103) );
  OA21x2_ASAP7_75t_R   g6425( .A1 (n6293), .A2 (n4754), .B (n3302), .Y (y3104) );
  AO21x1_ASAP7_75t_R   g6426( .A1 (n17), .A2 (x0), .B (x1), .Y (n6434) );
  AND2x2_ASAP7_75t_R   g6427( .A (n244), .B (n746), .Y (n6435) );
  INVx1_ASAP7_75t_R    g6428( .A (n6435), .Y (n6436) );
  AO21x1_ASAP7_75t_R   g6429( .A1 (n244), .A2 (n746), .B (x3), .Y (n6437) );
  OAI21x1_ASAP7_75t_R  g6430( .A1 (n17), .A2 (n6436), .B (n6437), .Y (n6438) );
  OA22x2_ASAP7_75t_R   g6431( .A1 (n6434), .A2 (n3033), .B1 (n6438), .B2 (n16), .Y (y3105) );
  AO221x2_ASAP7_75t_R  g6432( .A1 (x2), .A2 (n529), .B1 (n5177), .B2 (n4621), .C (n3294), .Y (y3106) );
  AO21x1_ASAP7_75t_R   g6433( .A1 (n369), .A2 (n388), .B (x2), .Y (n6441) );
  OA21x2_ASAP7_75t_R   g6434( .A1 (n3009), .A2 (n3237), .B (n6441), .Y (y3107) );
  INVx1_ASAP7_75t_R    g6435( .A (y1474), .Y (n6443) );
  NOR2x1_ASAP7_75t_R   g6436( .A (n6443), .B (y2071), .Y (y3108) );
  AND2x2_ASAP7_75t_R   g6437( .A (n3049), .B (n1720), .Y (y3109) );
  NAND2x1_ASAP7_75t_R  g6438( .A (n12), .B (n3376), .Y (n6446) );
  AND2x2_ASAP7_75t_R   g6439( .A (n3138), .B (n6446), .Y (y3110) );
  AND2x2_ASAP7_75t_R   g6440( .A (n3496), .B (n1077), .Y (y3111) );
  AO21x1_ASAP7_75t_R   g6441( .A1 (n455), .A2 (x2), .B (n5928), .Y (n6449) );
  OA21x2_ASAP7_75t_R   g6442( .A1 (n6234), .A2 (n5884), .B (n6449), .Y (y3112) );
  AND2x2_ASAP7_75t_R   g6443( .A (y168), .B (n3376), .Y (y3113) );
  AND2x2_ASAP7_75t_R   g6444( .A (n4014), .B (n22), .Y (n6452) );
  OA21x2_ASAP7_75t_R   g6445( .A1 (n6452), .A2 (n308), .B (n3882), .Y (y3114) );
  OR3x1_ASAP7_75t_R    g6446( .A (n999), .B (y2079), .C (n12), .Y (n6454) );
  INVx1_ASAP7_75t_R    g6447( .A (n6454), .Y (n6455) );
  AO21x1_ASAP7_75t_R   g6448( .A1 (n28), .A2 (n1208), .B (n6455), .Y (n6456) );
  XOR2x2_ASAP7_75t_R   g6449( .A (n6456), .B (x4), .Y (y3115) );
  OA21x2_ASAP7_75t_R   g6450( .A1 (n5250), .A2 (n15), .B (n4022), .Y (y3116) );
  AND3x1_ASAP7_75t_R   g6451( .A (n6272), .B (n72), .C (n5522), .Y (y3117) );
  OR3x1_ASAP7_75t_R    g6452( .A (n1158), .B (n291), .C (y2079), .Y (n6460) );
  AND2x2_ASAP7_75t_R   g6453( .A (n656), .B (n661), .Y (n6461) );
  AND2x2_ASAP7_75t_R   g6454( .A (n6460), .B (n6461), .Y (y3118) );
  OR3x1_ASAP7_75t_R    g6455( .A (n58), .B (x3), .C (x4), .Y (n6463) );
  AND2x2_ASAP7_75t_R   g6456( .A (n6463), .B (n5828), .Y (y3119) );
  OA21x2_ASAP7_75t_R   g6457( .A1 (n5250), .A2 (n15), .B (n3238), .Y (y3120) );
  AO21x1_ASAP7_75t_R   g6458( .A1 (y3852), .A2 (n22), .B (n3645), .Y (n6466) );
  OA21x2_ASAP7_75t_R   g6459( .A1 (n1112), .A2 (x3), .B (n6466), .Y (y3121) );
  AO21x1_ASAP7_75t_R   g6460( .A1 (n856), .A2 (n228), .B (y2393), .Y (y3122) );
  AND2x2_ASAP7_75t_R   g6461( .A (n366), .B (x2), .Y (n6469) );
  AO21x1_ASAP7_75t_R   g6462( .A1 (n388), .A2 (n45), .B (n6469), .Y (y3123) );
  OA33x2_ASAP7_75t_R   g6463( .A1 (n17), .A2 (y2079), .A3 (x2), .B1 (n3819), .B2 (n1158), .B3 (n1646), .Y (y3124) );
  OR3x1_ASAP7_75t_R    g6464( .A (n145), .B (n16), .C (n15), .Y (n6472) );
  AO21x1_ASAP7_75t_R   g6465( .A1 (n762), .A2 (n17), .B (n13), .Y (n6473) );
  AND2x2_ASAP7_75t_R   g6466( .A (n6472), .B (n6473), .Y (y3125) );
  NAND2x1_ASAP7_75t_R  g6467( .A (n4109), .B (n6326), .Y (y3126) );
  AND3x1_ASAP7_75t_R   g6468( .A (n1062), .B (n3024), .C (n556), .Y (n6476) );
  AO21x1_ASAP7_75t_R   g6469( .A1 (x4), .A2 (n3294), .B (n6476), .Y (y3128) );
  AND3x1_ASAP7_75t_R   g6470( .A (y3397), .B (n672), .C (n3000), .Y (y3129) );
  AND3x1_ASAP7_75t_R   g6471( .A (n1039), .B (n219), .C (y3293), .Y (y3130) );
  AND2x2_ASAP7_75t_R   g6472( .A (n455), .B (n72), .Y (n6480) );
  AND2x2_ASAP7_75t_R   g6473( .A (n3302), .B (n6480), .Y (y3131) );
  AO21x1_ASAP7_75t_R   g6474( .A1 (n455), .A2 (n72), .B (n163), .Y (n6482) );
  AND2x2_ASAP7_75t_R   g6475( .A (n3302), .B (n6482), .Y (y3133) );
  OR3x1_ASAP7_75t_R    g6476( .A (n5307), .B (y2079), .C (y863), .Y (y3135) );
  AO21x1_ASAP7_75t_R   g6477( .A1 (n1564), .A2 (n63), .B (n363), .Y (y3136) );
  AND2x2_ASAP7_75t_R   g6478( .A (n3302), .B (n6351), .Y (y3137) );
  AO32x1_ASAP7_75t_R   g6479( .A1 (n72), .A2 (n3585), .A3 (n4495), .B1 (n4109), .B2 (n6287), .Y (n6487) );
  INVx1_ASAP7_75t_R    g6480( .A (n6487), .Y (y3138) );
  NAND2x1_ASAP7_75t_R  g6481( .A (n15), .B (n3457), .Y (n6489) );
  AND2x2_ASAP7_75t_R   g6482( .A (n3302), .B (n6489), .Y (y3139) );
  AND3x1_ASAP7_75t_R   g6483( .A (n2296), .B (n2141), .C (n244), .Y (y3140) );
  NOR2x1_ASAP7_75t_R   g6484( .A (n15), .B (n3218), .Y (n6492) );
  AO21x1_ASAP7_75t_R   g6485( .A1 (x5), .A2 (n3310), .B (n6492), .Y (y3141) );
  AND2x2_ASAP7_75t_R   g6486( .A (y3274), .B (n3577), .Y (y3142) );
  NAND2x1_ASAP7_75t_R  g6487( .A (n292), .B (n125), .Y (n6495) );
  AND2x2_ASAP7_75t_R   g6488( .A (n6495), .B (n4362), .Y (y3144) );
  AO21x1_ASAP7_75t_R   g6489( .A1 (n1158), .A2 (n97), .B (n3819), .Y (n6497) );
  AO21x1_ASAP7_75t_R   g6490( .A1 (n15), .A2 (n17), .B (n6497), .Y (y3145) );
  OAI21x1_ASAP7_75t_R  g6491( .A1 (n81), .A2 (n5446), .B (n3448), .Y (y3146) );
  INVx1_ASAP7_75t_R    g6492( .A (n4151), .Y (n6500) );
  OR3x1_ASAP7_75t_R    g6493( .A (n5427), .B (n1269), .C (n6500), .Y (y3147) );
  AND2x2_ASAP7_75t_R   g6494( .A (n3790), .B (n3805), .Y (y3148) );
  AO21x1_ASAP7_75t_R   g6495( .A1 (n366), .A2 (n5090), .B (n3294), .Y (y3149) );
  AND2x2_ASAP7_75t_R   g6496( .A (n28), .B (n3469), .Y (n6504) );
  OA21x2_ASAP7_75t_R   g6497( .A1 (n6504), .A2 (n4216), .B (y3340), .Y (y3150) );
  OA21x2_ASAP7_75t_R   g6498( .A1 (x5), .A2 (n3471), .B (y3171), .Y (y3151) );
  AO21x1_ASAP7_75t_R   g6499( .A1 (n3568), .A2 (x3), .B (n4502), .Y (y3169) );
  AND2x2_ASAP7_75t_R   g6500( .A (y3169), .B (n5507), .Y (y3152) );
  AND2x2_ASAP7_75t_R   g6501( .A (y3169), .B (n4504), .Y (y3153) );
  OR3x1_ASAP7_75t_R    g6502( .A (n628), .B (n638), .C (x0), .Y (y3154) );
  AO21x1_ASAP7_75t_R   g6503( .A1 (n22), .A2 (x5), .B (y863), .Y (n6511) );
  AO21x1_ASAP7_75t_R   g6504( .A1 (y2079), .A2 (n1707), .B (n6511), .Y (y3155) );
  OA21x2_ASAP7_75t_R   g6505( .A1 (n403), .A2 (n4022), .B (n5879), .Y (y3156) );
  OA21x2_ASAP7_75t_R   g6506( .A1 (n1337), .A2 (n5905), .B (n1440), .Y (y3157) );
  NAND2x1_ASAP7_75t_R  g6507( .A (n1166), .B (n1747), .Y (n6515) );
  AND2x2_ASAP7_75t_R   g6508( .A (n6515), .B (y1281), .Y (y3158) );
  AND2x2_ASAP7_75t_R   g6509( .A (n366), .B (n3143), .Y (n6517) );
  AO21x1_ASAP7_75t_R   g6510( .A1 (n388), .A2 (n45), .B (n6517), .Y (y3159) );
  AND3x1_ASAP7_75t_R   g6511( .A (n4469), .B (n5520), .C (y1359), .Y (y3161) );
  OR3x1_ASAP7_75t_R    g6512( .A (n529), .B (n17), .C (n756), .Y (n6520) );
  OA21x2_ASAP7_75t_R   g6513( .A1 (n529), .A2 (n4495), .B (n6520), .Y (y3162) );
  OR3x1_ASAP7_75t_R    g6514( .A (n143), .B (y2079), .C (n22), .Y (n6522) );
  AND2x2_ASAP7_75t_R   g6515( .A (n453), .B (n6522), .Y (y3163) );
  INVx1_ASAP7_75t_R    g6516( .A (n6045), .Y (n6524) );
  AND2x2_ASAP7_75t_R   g6517( .A (n5127), .B (y2079), .Y (n6525) );
  AO21x1_ASAP7_75t_R   g6518( .A1 (n3685), .A2 (n6524), .B (n6525), .Y (y3164) );
  AND2x2_ASAP7_75t_R   g6519( .A (n1064), .B (n6522), .Y (y3165) );
  NAND2x1_ASAP7_75t_R  g6520( .A (n17), .B (n3466), .Y (n6528) );
  OA21x2_ASAP7_75t_R   g6521( .A1 (n2843), .A2 (n17), .B (n6528), .Y (y3166) );
  AO21x1_ASAP7_75t_R   g6522( .A1 (n17), .A2 (n757), .B (n2990), .Y (y3167) );
  AO32x1_ASAP7_75t_R   g6523( .A1 (x5), .A2 (n72), .A3 (n4495), .B1 (y2079), .B2 (n5181), .Y (y3168) );
  NOR2x1_ASAP7_75t_R   g6524( .A (y2498), .B (n3439), .Y (y3170) );
  AO21x1_ASAP7_75t_R   g6525( .A1 (x0), .A2 (n556), .B (n4679), .Y (y3172) );
  INVx1_ASAP7_75t_R    g6526( .A (n4325), .Y (n6534) );
  NOR2x1_ASAP7_75t_R   g6527( .A (n6534), .B (n4736), .Y (n6535) );
  AO21x1_ASAP7_75t_R   g6528( .A1 (n360), .A2 (y2079), .B (n3359), .Y (n6536) );
  OA21x2_ASAP7_75t_R   g6529( .A1 (n6535), .A2 (x2), .B (n6536), .Y (y3173) );
  AO32x1_ASAP7_75t_R   g6530( .A1 (n3524), .A2 (x5), .A3 (n3000), .B1 (n3585), .B2 (n3705), .Y (y3174) );
  OR3x1_ASAP7_75t_R    g6531( .A (y3758), .B (n15), .C (n1158), .Y (n6539) );
  OA21x2_ASAP7_75t_R   g6532( .A1 (x2), .A2 (n389), .B (n6539), .Y (y3175) );
  OA21x2_ASAP7_75t_R   g6533( .A1 (n389), .A2 (x2), .B (n4341), .Y (y3177) );
  AO21x1_ASAP7_75t_R   g6534( .A1 (y3293), .A2 (x0), .B (n410), .Y (n6542) );
  OA21x2_ASAP7_75t_R   g6535( .A1 (x1), .A2 (n6542), .B (n935), .Y (y3178) );
  OA21x2_ASAP7_75t_R   g6536( .A1 (n1158), .A2 (n5001), .B (y3276), .Y (y3179) );
  AND3x1_ASAP7_75t_R   g6537( .A (n1062), .B (n3823), .C (y3293), .Y (n6545) );
  AO21x1_ASAP7_75t_R   g6538( .A1 (x5), .A2 (n3263), .B (n6545), .Y (y3180) );
  AO32x1_ASAP7_75t_R   g6539( .A1 (n360), .A2 (n5055), .A3 (n290), .B1 (n4225), .B2 (n4681), .Y (y3181) );
  INVx1_ASAP7_75t_R    g6540( .A (n2665), .Y (n6548) );
  OA21x2_ASAP7_75t_R   g6541( .A1 (n6548), .A2 (x4), .B (n496), .Y (y3182) );
  AO21x1_ASAP7_75t_R   g6542( .A1 (n128), .A2 (n481), .B (y1206), .Y (y3183) );
  INVx1_ASAP7_75t_R    g6543( .A (n4366), .Y (n6551) );
  AND2x2_ASAP7_75t_R   g6544( .A (y3276), .B (n6551), .Y (y3184) );
  NOR2x1_ASAP7_75t_R   g6545( .A (n4340), .B (n5482), .Y (y3185) );
  OA22x2_ASAP7_75t_R   g6546( .A1 (n4695), .A2 (n4788), .B1 (n3278), .B2 (n22), .Y (y3186) );
  AO21x1_ASAP7_75t_R   g6547( .A1 (n740), .A2 (n4621), .B (n4841), .Y (y3187) );
  AO21x1_ASAP7_75t_R   g6548( .A1 (n316), .A2 (n22), .B (n3237), .Y (n6556) );
  OA21x2_ASAP7_75t_R   g6549( .A1 (n4586), .A2 (n3377), .B (n6556), .Y (y3188) );
  OR3x1_ASAP7_75t_R    g6550( .A (n81), .B (x1), .C (x0), .Y (n6558) );
  AND2x2_ASAP7_75t_R   g6551( .A (n1697), .B (n6558), .Y (y3189) );
  NAND2x1_ASAP7_75t_R  g6552( .A (n15), .B (n5730), .Y (n6560) );
  AND2x2_ASAP7_75t_R   g6553( .A (n6539), .B (n6560), .Y (y3190) );
  AND2x2_ASAP7_75t_R   g6554( .A (n4341), .B (n3377), .Y (y3191) );
  AND3x1_ASAP7_75t_R   g6555( .A (n221), .B (n17), .C (n15), .Y (n6563) );
  AO21x1_ASAP7_75t_R   g6556( .A1 (n2432), .A2 (n2271), .B (n6563), .Y (y3192) );
  AO21x1_ASAP7_75t_R   g6557( .A1 (n6404), .A2 (n5090), .B (n3263), .Y (y3193) );
  INVx1_ASAP7_75t_R    g6558( .A (n2600), .Y (n6566) );
  AND2x2_ASAP7_75t_R   g6559( .A (y3134), .B (n6566), .Y (y3194) );
  OA21x2_ASAP7_75t_R   g6560( .A1 (n518), .A2 (n4238), .B (y3397), .Y (y3195) );
  AND3x1_ASAP7_75t_R   g6561( .A (n316), .B (n319), .C (n22), .Y (n6569) );
  OR3x1_ASAP7_75t_R    g6562( .A (n321), .B (n6569), .C (n323), .Y (y3196) );
  AO221x2_ASAP7_75t_R  g6563( .A1 (n45), .A2 (n1545), .B1 (n144), .B2 (n218), .C (n2588), .Y (y3197) );
  NOR2x1_ASAP7_75t_R   g6564( .A (n5801), .B (n6291), .Y (n6572) );
  OR3x1_ASAP7_75t_R    g6565( .A (n6572), .B (n3443), .C (n3279), .Y (y3199) );
  AO21x1_ASAP7_75t_R   g6566( .A1 (y9), .A2 (n29), .B (n4808), .Y (y3200) );
  OA22x2_ASAP7_75t_R   g6567( .A1 (n5323), .A2 (n4695), .B1 (n3294), .B2 (n4903), .Y (y3201) );
  NAND2x1_ASAP7_75t_R  g6568( .A (x0), .B (n705), .Y (n6576) );
  AND2x2_ASAP7_75t_R   g6569( .A (n6576), .B (n707), .Y (y3202) );
  OA21x2_ASAP7_75t_R   g6570( .A1 (n403), .A2 (n4528), .B (n5879), .Y (y3203) );
  INVx1_ASAP7_75t_R    g6571( .A (n370), .Y (n6579) );
  AO21x1_ASAP7_75t_R   g6572( .A1 (n6579), .A2 (n3023), .B (n3568), .Y (y3204) );
  AO21x1_ASAP7_75t_R   g6573( .A1 (n5085), .A2 (n3377), .B (n628), .Y (y3205) );
  NAND2x1_ASAP7_75t_R  g6574( .A (x5), .B (n3267), .Y (n6582) );
  AO21x1_ASAP7_75t_R   g6575( .A1 (n6582), .A2 (n299), .B (n3080), .Y (y3206) );
  AO21x1_ASAP7_75t_R   g6576( .A1 (y2079), .A2 (x0), .B (n43), .Y (n6584) );
  AO21x1_ASAP7_75t_R   g6577( .A1 (n6584), .A2 (x2), .B (n1778), .Y (y3207) );
  AO21x1_ASAP7_75t_R   g6578( .A1 (n1492), .A2 (n4625), .B (n2193), .Y (n6586) );
  AO21x1_ASAP7_75t_R   g6579( .A1 (n12), .A2 (n15), .B (n6586), .Y (y3208) );
  AND2x2_ASAP7_75t_R   g6580( .A (n4111), .B (n5843), .Y (y3209) );
  OA21x2_ASAP7_75t_R   g6581( .A1 (x0), .A2 (n552), .B (n5114), .Y (y3210) );
  OR3x1_ASAP7_75t_R    g6582( .A (n3296), .B (n4621), .C (n628), .Y (y3211) );
  AND2x2_ASAP7_75t_R   g6583( .A (n290), .B (n4117), .Y (n6591) );
  INVx1_ASAP7_75t_R    g6584( .A (n6591), .Y (n6592) );
  AO21x1_ASAP7_75t_R   g6585( .A1 (n1851), .A2 (n17), .B (n366), .Y (n6593) );
  INVx1_ASAP7_75t_R    g6586( .A (n6593), .Y (n6594) );
  AO21x1_ASAP7_75t_R   g6587( .A1 (y2079), .A2 (n6592), .B (n6594), .Y (n6595) );
  NAND2x1_ASAP7_75t_R  g6588( .A (n328), .B (n6595), .Y (y3212) );
  AO21x1_ASAP7_75t_R   g6589( .A1 (n989), .A2 (x2), .B (n128), .Y (y3213) );
  OA21x2_ASAP7_75t_R   g6590( .A1 (n5654), .A2 (n22), .B (n4695), .Y (y3214) );
  AND2x2_ASAP7_75t_R   g6591( .A (y117), .B (n419), .Y (y3215) );
  OA21x2_ASAP7_75t_R   g6592( .A1 (n3443), .A2 (n5707), .B (n4056), .Y (y3216) );
  AO21x1_ASAP7_75t_R   g6593( .A1 (y2079), .A2 (n4647), .B (n3992), .Y (n6601) );
  AO21x1_ASAP7_75t_R   g6594( .A1 (x5), .A2 (n4648), .B (n6601), .Y (y3217) );
  OA21x2_ASAP7_75t_R   g6595( .A1 (n22), .A2 (n5654), .B (n4904), .Y (y3218) );
  INVx1_ASAP7_75t_R    g6596( .A (n3694), .Y (n6604) );
  AND2x2_ASAP7_75t_R   g6597( .A (y2958), .B (n6604), .Y (y3219) );
  AO21x1_ASAP7_75t_R   g6598( .A1 (n22), .A2 (x2), .B (y2079), .Y (n6606) );
  INVx1_ASAP7_75t_R    g6599( .A (n6606), .Y (n6607) );
  AOI22x1_ASAP7_75t_R  g6600( .A1 (n4518), .A2 (n3474), .B1 (n6607), .B2 (n290), .Y (y3220) );
  INVx1_ASAP7_75t_R    g6601( .A (n2994), .Y (n6609) );
  AO21x1_ASAP7_75t_R   g6602( .A1 (n22), .A2 (x3), .B (n2994), .Y (n6610) );
  AO32x1_ASAP7_75t_R   g6603( .A1 (n360), .A2 (n6609), .A3 (y2079), .B1 (x5), .B2 (n6610), .Y (y3221) );
  NOR2x1_ASAP7_75t_R   g6604( .A (n316), .B (n3567), .Y (n6612) );
  INVx1_ASAP7_75t_R    g6605( .A (n6612), .Y (n6613) );
  AND2x2_ASAP7_75t_R   g6606( .A (n6613), .B (y2958), .Y (y3222) );
  AO21x1_ASAP7_75t_R   g6607( .A1 (n368), .A2 (x4), .B (x2), .Y (n6615) );
  OA21x2_ASAP7_75t_R   g6608( .A1 (n3474), .A2 (n4495), .B (n6615), .Y (y3223) );
  OR3x1_ASAP7_75t_R    g6609( .A (n798), .B (y2079), .C (n61), .Y (n6617) );
  AND2x2_ASAP7_75t_R   g6610( .A (n6617), .B (n6576), .Y (y3224) );
  OA21x2_ASAP7_75t_R   g6611( .A1 (n4361), .A2 (n45), .B (n3000), .Y (y3225) );
  AND3x1_ASAP7_75t_R   g6612( .A (n656), .B (n2984), .C (n5843), .Y (y3226) );
  AO21x1_ASAP7_75t_R   g6613( .A1 (n672), .A2 (n4640), .B (n3272), .Y (y3227) );
  AO21x1_ASAP7_75t_R   g6614( .A1 (n5654), .A2 (x4), .B (n3568), .Y (y3228) );
  OA22x2_ASAP7_75t_R   g6615( .A1 (n701), .A2 (n2503), .B1 (n2508), .B2 (n16), .Y (y3229) );
  AO21x1_ASAP7_75t_R   g6616( .A1 (n22), .A2 (x2), .B (n3443), .Y (n6624) );
  AO21x1_ASAP7_75t_R   g6617( .A1 (n45), .A2 (n28), .B (n6624), .Y (y3230) );
  OR3x1_ASAP7_75t_R    g6618( .A (n3272), .B (n3279), .C (n628), .Y (y3231) );
  AO21x1_ASAP7_75t_R   g6619( .A1 (n4083), .A2 (n556), .B (n1137), .Y (y3232) );
  OA21x2_ASAP7_75t_R   g6620( .A1 (n291), .A2 (n6606), .B (n4536), .Y (y3233) );
  OA21x2_ASAP7_75t_R   g6621( .A1 (n6579), .A2 (n4273), .B (y3397), .Y (y3235) );
  AND3x1_ASAP7_75t_R   g6622( .A (n4016), .B (n3882), .C (n299), .Y (y3236) );
  OR3x1_ASAP7_75t_R    g6623( .A (n1000), .B (n231), .C (x0), .Y (y3237) );
  OA21x2_ASAP7_75t_R   g6624( .A1 (n1277), .A2 (n3636), .B (n6556), .Y (y3238) );
  OA21x2_ASAP7_75t_R   g6625( .A1 (n5633), .A2 (n3414), .B (n3648), .Y (y3239) );
  INVx1_ASAP7_75t_R    g6626( .A (n3263), .Y (n6634) );
  AO21x1_ASAP7_75t_R   g6627( .A1 (n3777), .A2 (x2), .B (n3263), .Y (n6635) );
  AO32x1_ASAP7_75t_R   g6628( .A1 (n6634), .A2 (n3550), .A3 (y2079), .B1 (x5), .B2 (n6635), .Y (y3240) );
  NAND2x1_ASAP7_75t_R  g6629( .A (n844), .B (n3840), .Y (y3241) );
  AND3x1_ASAP7_75t_R   g6630( .A (y3397), .B (n5148), .C (n3000), .Y (y3242) );
  OA21x2_ASAP7_75t_R   g6631( .A1 (n2511), .A2 (n1209), .B (n1490), .Y (y3243) );
  AND2x2_ASAP7_75t_R   g6632( .A (n378), .B (y2079), .Y (y3244) );
  AO21x1_ASAP7_75t_R   g6633( .A1 (n382), .A2 (y3852), .B (y2196), .Y (y3245) );
  AO21x1_ASAP7_75t_R   g6634( .A1 (n45), .A2 (n28), .B (n4640), .Y (y3267) );
  AO21x1_ASAP7_75t_R   g6635( .A1 (n3469), .A2 (n3567), .B (n672), .Y (n6643) );
  AND2x2_ASAP7_75t_R   g6636( .A (y3267), .B (n6643), .Y (y3246) );
  AO21x1_ASAP7_75t_R   g6637( .A1 (x5), .A2 (n537), .B (n418), .Y (n6645) );
  AO21x1_ASAP7_75t_R   g6638( .A1 (n17), .A2 (n6645), .B (n3062), .Y (y3247) );
  AO21x1_ASAP7_75t_R   g6639( .A1 (n3023), .A2 (n5507), .B (n22), .Y (n6647) );
  OA21x2_ASAP7_75t_R   g6640( .A1 (n671), .A2 (n3000), .B (n6647), .Y (y3248) );
  NOR2x1_ASAP7_75t_R   g6641( .A (n12), .B (n5968), .Y (y3249) );
  AND2x2_ASAP7_75t_R   g6642( .A (y2708), .B (n4737), .Y (y3250) );
  OR3x1_ASAP7_75t_R    g6643( .A (n291), .B (n5108), .C (y2079), .Y (n6651) );
  AO32x1_ASAP7_75t_R   g6644( .A1 (n290), .A2 (n3207), .A3 (n15), .B1 (x2), .B2 (n6651), .Y (y3251) );
  AO32x1_ASAP7_75t_R   g6645( .A1 (n3028), .A2 (n3377), .A3 (x5), .B1 (y2079), .B2 (n4924), .Y (y3252) );
  NAND2x1_ASAP7_75t_R  g6646( .A (n3905), .B (n3866), .Y (n6654) );
  AO21x1_ASAP7_75t_R   g6647( .A1 (x4), .A2 (n3294), .B (n6654), .Y (y3253) );
  AND2x2_ASAP7_75t_R   g6648( .A (y1474), .B (n6604), .Y (y3254) );
  AND2x2_ASAP7_75t_R   g6649( .A (n3023), .B (x4), .Y (n6657) );
  AO21x1_ASAP7_75t_R   g6650( .A1 (n22), .A2 (n4273), .B (n6657), .Y (y3255) );
  INVx1_ASAP7_75t_R    g6651( .A (n3023), .Y (n6659) );
  OA21x2_ASAP7_75t_R   g6652( .A1 (n6659), .A2 (n4844), .B (y1474), .Y (y3256) );
  OA21x2_ASAP7_75t_R   g6653( .A1 (n3611), .A2 (n22), .B (n4109), .Y (y3257) );
  AO21x1_ASAP7_75t_R   g6654( .A1 (n3023), .A2 (n4844), .B (n4042), .Y (y3258) );
  OA21x2_ASAP7_75t_R   g6655( .A1 (n2321), .A2 (x1), .B (n733), .Y (y3259) );
  NOR2x1_ASAP7_75t_R   g6656( .A (n3694), .B (n6607), .Y (n6664) );
  AO21x1_ASAP7_75t_R   g6657( .A1 (n17), .A2 (n3183), .B (n6664), .Y (y3260) );
  AO21x1_ASAP7_75t_R   g6658( .A1 (x4), .A2 (x5), .B (x0), .Y (n6666) );
  INVx1_ASAP7_75t_R    g6659( .A (n6666), .Y (n6667) );
  AO21x1_ASAP7_75t_R   g6660( .A1 (n360), .A2 (n6667), .B (n3269), .Y (y3261) );
  OA21x2_ASAP7_75t_R   g6661( .A1 (x4), .A2 (n3556), .B (y3397), .Y (y3263) );
  AND3x1_ASAP7_75t_R   g6662( .A (n45), .B (y2079), .C (n22), .Y (y3264) );
  AO21x1_ASAP7_75t_R   g6663( .A1 (n45), .A2 (n28), .B (n4995), .Y (y3265) );
  AND2x2_ASAP7_75t_R   g6664( .A (y3397), .B (n3000), .Y (y3266) );
  AND2x2_ASAP7_75t_R   g6665( .A (y3245), .B (n5493), .Y (y3268) );
  OA21x2_ASAP7_75t_R   g6666( .A1 (n529), .A2 (n3341), .B (n642), .Y (y3270) );
  INVx1_ASAP7_75t_R    g6667( .A (n3550), .Y (n6675) );
  AO21x1_ASAP7_75t_R   g6668( .A1 (n3023), .A2 (n3123), .B (n6675), .Y (y3271) );
  AO21x1_ASAP7_75t_R   g6669( .A1 (n1894), .A2 (x0), .B (n1896), .Y (y3272) );
  NAND2x1_ASAP7_75t_R  g6670( .A (n3526), .B (n3524), .Y (n6678) );
  AO21x1_ASAP7_75t_R   g6671( .A1 (n3524), .A2 (n3526), .B (y2079), .Y (n6679) );
  OA21x2_ASAP7_75t_R   g6672( .A1 (n6678), .A2 (n1265), .B (n6679), .Y (y3273) );
  AO32x1_ASAP7_75t_R   g6673( .A1 (y103), .A2 (n934), .A3 (n3014), .B1 (x3), .B2 (y1378), .Y (y3275) );
  AND2x2_ASAP7_75t_R   g6674( .A (n221), .B (n17), .Y (n6682) );
  OA21x2_ASAP7_75t_R   g6675( .A1 (n2583), .A2 (n243), .B (n1480), .Y (n6683) );
  AO21x1_ASAP7_75t_R   g6676( .A1 (n6682), .A2 (n15), .B (n6683), .Y (y3277) );
  AO32x1_ASAP7_75t_R   g6677( .A1 (n3377), .A2 (x5), .A3 (n3028), .B1 (n5385), .B2 (n6634), .Y (y3278) );
  AND3x1_ASAP7_75t_R   g6678( .A (n3013), .B (n72), .C (n419), .Y (y3279) );
  AND2x2_ASAP7_75t_R   g6679( .A (n1590), .B (n2848), .Y (n6687) );
  NOR2x1_ASAP7_75t_R   g6680( .A (n2718), .B (n6687), .Y (y3280) );
  OR3x1_ASAP7_75t_R    g6681( .A (n403), .B (y2079), .C (n12), .Y (n6689) );
  INVx1_ASAP7_75t_R    g6682( .A (n6689), .Y (n6690) );
  OR3x1_ASAP7_75t_R    g6683( .A (n6690), .B (n676), .C (n337), .Y (y3281) );
  AO21x1_ASAP7_75t_R   g6684( .A1 (y3758), .A2 (x2), .B (n6218), .Y (y3282) );
  AO21x1_ASAP7_75t_R   g6685( .A1 (n15), .A2 (n401), .B (n163), .Y (n6693) );
  INVx1_ASAP7_75t_R    g6686( .A (n6693), .Y (n6694) );
  AO21x1_ASAP7_75t_R   g6687( .A1 (y2079), .A2 (n6694), .B (n4114), .Y (y3283) );
  INVx1_ASAP7_75t_R    g6688( .A (n3132), .Y (n6696) );
  AO21x1_ASAP7_75t_R   g6689( .A1 (n6696), .A2 (n6010), .B (n4243), .Y (y3284) );
  AND3x1_ASAP7_75t_R   g6690( .A (n2999), .B (y2079), .C (x3), .Y (n6698) );
  AO21x1_ASAP7_75t_R   g6691( .A1 (n6480), .A2 (n4341), .B (n6698), .Y (y3285) );
  AND2x2_ASAP7_75t_R   g6692( .A (n4548), .B (n3459), .Y (y3286) );
  NAND2x1_ASAP7_75t_R  g6693( .A (n292), .B (n319), .Y (n6701) );
  XOR2x2_ASAP7_75t_R   g6694( .A (n6701), .B (n5227), .Y (y3287) );
  NAND2x1_ASAP7_75t_R  g6695( .A (n15), .B (n391), .Y (n6703) );
  OA21x2_ASAP7_75t_R   g6696( .A1 (n6703), .A2 (n959), .B (n6536), .Y (y3288) );
  AND2x2_ASAP7_75t_R   g6697( .A (n6536), .B (n3825), .Y (y3289) );
  AND3x1_ASAP7_75t_R   g6698( .A (n3013), .B (n72), .C (n3832), .Y (y3290) );
  AND2x2_ASAP7_75t_R   g6699( .A (y1903), .B (n3977), .Y (y3291) );
  AND2x2_ASAP7_75t_R   g6700( .A (n6539), .B (n72), .Y (y3292) );
  AO21x1_ASAP7_75t_R   g6701( .A1 (n369), .A2 (n299), .B (n914), .Y (n6709) );
  OA21x2_ASAP7_75t_R   g6702( .A1 (n407), .A2 (n409), .B (n6709), .Y (y3294) );
  OA33x2_ASAP7_75t_R   g6703( .A1 (x5), .A2 (n403), .A3 (n3375), .B1 (y2079), .B2 (n3263), .B3 (n5427), .Y (y3295) );
  AO21x1_ASAP7_75t_R   g6704( .A1 (n6480), .A2 (n4341), .B (n4586), .Y (y3296) );
  AND2x2_ASAP7_75t_R   g6705( .A (y3293), .B (n3823), .Y (n6713) );
  OA21x2_ASAP7_75t_R   g6706( .A1 (n45), .A2 (n6713), .B (n4031), .Y (y3297) );
  AND2x2_ASAP7_75t_R   g6707( .A (n5090), .B (n366), .Y (n6715) );
  AO21x1_ASAP7_75t_R   g6708( .A1 (x4), .A2 (n3294), .B (n6715), .Y (y3298) );
  AND2x2_ASAP7_75t_R   g6709( .A (y2610), .B (n455), .Y (y3299) );
  OR3x1_ASAP7_75t_R    g6710( .A (n3443), .B (n3279), .C (n45), .Y (y3300) );
  AO21x1_ASAP7_75t_R   g6711( .A1 (n3366), .A2 (y2079), .B (n143), .Y (n6719) );
  AO21x1_ASAP7_75t_R   g6712( .A1 (n481), .A2 (n527), .B (n6719), .Y (y3301) );
  OA211x2_ASAP7_75t_R  g6713( .A1 (n5072), .A2 (n914), .B (n3884), .C (n5342), .Y (y3302) );
  AO32x1_ASAP7_75t_R   g6714( .A1 (n285), .A2 (n287), .A3 (n15), .B1 (x2), .B2 (y3808), .Y (y3303) );
  OR3x1_ASAP7_75t_R    g6715( .A (n4042), .B (n3443), .C (n45), .Y (y3304) );
  AND2x2_ASAP7_75t_R   g6716( .A (y3397), .B (n5756), .Y (y3306) );
  AND2x2_ASAP7_75t_R   g6717( .A (y2432), .B (n475), .Y (y3307) );
  XOR2x2_ASAP7_75t_R   g6718( .A (n6326), .B (n3024), .Y (y3308) );
  AND3x1_ASAP7_75t_R   g6719( .A (n360), .B (n290), .C (n15), .Y (n6727) );
  AO21x1_ASAP7_75t_R   g6720( .A1 (n5828), .A2 (x2), .B (n6727), .Y (y3309) );
  INVx1_ASAP7_75t_R    g6721( .A (n1296), .Y (n6729) );
  AO21x1_ASAP7_75t_R   g6722( .A1 (n12), .A2 (x2), .B (n143), .Y (n6730) );
  NAND2x1_ASAP7_75t_R  g6723( .A (x2), .B (n1253), .Y (n6731) );
  OA21x2_ASAP7_75t_R   g6724( .A1 (n6729), .A2 (n6730), .B (n6731), .Y (y3310) );
  INVx1_ASAP7_75t_R    g6725( .A (n5476), .Y (n6733) );
  OA21x2_ASAP7_75t_R   g6726( .A1 (n3750), .A2 (n6733), .B (y2610), .Y (y3311) );
  AND2x2_ASAP7_75t_R   g6727( .A (n6613), .B (y2610), .Y (y3312) );
  AO21x1_ASAP7_75t_R   g6728( .A1 (n4640), .A2 (n5179), .B (n3294), .Y (y3313) );
  AO21x1_ASAP7_75t_R   g6729( .A1 (n436), .A2 (x0), .B (n3423), .Y (n6737) );
  AO32x1_ASAP7_75t_R   g6730( .A1 (n2008), .A2 (n3424), .A3 (n29), .B1 (y2079), .B2 (n6737), .Y (y3314) );
  INVx1_ASAP7_75t_R    g6731( .A (n4403), .Y (n6739) );
  AND2x2_ASAP7_75t_R   g6732( .A (n6739), .B (y2085), .Y (y3315) );
  AO21x1_ASAP7_75t_R   g6733( .A1 (n4640), .A2 (n672), .B (n45), .Y (y3316) );
  AO21x1_ASAP7_75t_R   g6734( .A1 (n455), .A2 (n5654), .B (n3568), .Y (y3317) );
  OR3x1_ASAP7_75t_R    g6735( .A (n4554), .B (n3009), .C (n315), .Y (y3318) );
  OR3x1_ASAP7_75t_R    g6736( .A (n5534), .B (n306), .C (y2196), .Y (y3319) );
  AO21x1_ASAP7_75t_R   g6737( .A1 (n527), .A2 (y2079), .B (n143), .Y (y3320) );
  NOR2x1_ASAP7_75t_R   g6738( .A (n12), .B (n103), .Y (n6746) );
  INVx1_ASAP7_75t_R    g6739( .A (n1146), .Y (n6747) );
  OA21x2_ASAP7_75t_R   g6740( .A1 (n2889), .A2 (n6746), .B (n6747), .Y (n6748) );
  NOR2x1_ASAP7_75t_R   g6741( .A (n1032), .B (n6748), .Y (y3321) );
  AO21x1_ASAP7_75t_R   g6742( .A1 (n1062), .A2 (n529), .B (n3751), .Y (y3322) );
  OA21x2_ASAP7_75t_R   g6743( .A1 (x5), .A2 (n3471), .B (y1474), .Y (y3323) );
  NOR2x1_ASAP7_75t_R   g6744( .A (n481), .B (n3723), .Y (y3324) );
  AO21x1_ASAP7_75t_R   g6745( .A1 (n6604), .A2 (n6606), .B (n3263), .Y (y3325) );
  OR3x1_ASAP7_75t_R    g6746( .A (n4831), .B (n3263), .C (y2466), .Y (y3326) );
  AO21x1_ASAP7_75t_R   g6747( .A1 (n6634), .A2 (n5385), .B (n3751), .Y (y3327) );
  AO21x1_ASAP7_75t_R   g6748( .A1 (n1062), .A2 (n5859), .B (n3751), .Y (y3328) );
  AND3x1_ASAP7_75t_R   g6749( .A (n1863), .B (y195), .C (n466), .Y (y3329) );
  NOR2x1_ASAP7_75t_R   g6750( .A (n6443), .B (y2457), .Y (y3330) );
  AO21x1_ASAP7_75t_R   g6751( .A1 (n1046), .A2 (x0), .B (n3974), .Y (y3331) );
  AO32x1_ASAP7_75t_R   g6752( .A1 (n672), .A2 (n72), .A3 (n3028), .B1 (n1062), .B2 (n529), .Y (y3332) );
  OA21x2_ASAP7_75t_R   g6753( .A1 (x1), .A2 (n2060), .B (n1345), .Y (y3333) );
  AND2x2_ASAP7_75t_R   g6754( .A (x2), .B (x0), .Y (n6762) );
  AO21x1_ASAP7_75t_R   g6755( .A1 (n16), .A2 (n15), .B (n6762), .Y (n6763) );
  AO21x1_ASAP7_75t_R   g6756( .A1 (n16), .A2 (x0), .B (n17), .Y (n6764) );
  INVx1_ASAP7_75t_R    g6757( .A (n6764), .Y (n6765) );
  AO21x1_ASAP7_75t_R   g6758( .A1 (y863), .A2 (x2), .B (x3), .Y (n6766) );
  INVx1_ASAP7_75t_R    g6759( .A (n6766), .Y (n6767) );
  AO21x1_ASAP7_75t_R   g6760( .A1 (n6763), .A2 (n6765), .B (n6767), .Y (y3334) );
  OR3x1_ASAP7_75t_R    g6761( .A (n3867), .B (n3568), .C (n3294), .Y (y3335) );
  AND2x2_ASAP7_75t_R   g6762( .A (n6404), .B (n4109), .Y (y3336) );
  AO21x1_ASAP7_75t_R   g6763( .A1 (y2079), .A2 (n3629), .B (n3751), .Y (y3337) );
  OR3x1_ASAP7_75t_R    g6764( .A (n5539), .B (n4781), .C (n628), .Y (y3338) );
  AO21x1_ASAP7_75t_R   g6765( .A1 (y2079), .A2 (x4), .B (n3751), .Y (y3339) );
  OR3x1_ASAP7_75t_R    g6766( .A (n145), .B (n22), .C (y2079), .Y (n6774) );
  INVx1_ASAP7_75t_R    g6767( .A (n4305), .Y (n6775) );
  AO21x1_ASAP7_75t_R   g6768( .A1 (n6775), .A2 (x5), .B (y2498), .Y (n6776) );
  AO32x1_ASAP7_75t_R   g6769( .A1 (n1370), .A2 (n6774), .A3 (x3), .B1 (n17), .B2 (n6776), .Y (y3341) );
  AO21x1_ASAP7_75t_R   g6770( .A1 (n17), .A2 (x2), .B (x5), .Y (n6778) );
  INVx1_ASAP7_75t_R    g6771( .A (n6778), .Y (n6779) );
  OR3x1_ASAP7_75t_R    g6772( .A (n1158), .B (n291), .C (n6779), .Y (y3342) );
  OA21x2_ASAP7_75t_R   g6773( .A1 (n3384), .A2 (n3085), .B (n3327), .Y (y3343) );
  INVx1_ASAP7_75t_R    g6774( .A (n4371), .Y (n6782) );
  OA21x2_ASAP7_75t_R   g6775( .A1 (n6782), .A2 (n2989), .B (n1062), .Y (n6783) );
  AO21x1_ASAP7_75t_R   g6776( .A1 (n3705), .A2 (n4371), .B (x5), .Y (n6784) );
  OA21x2_ASAP7_75t_R   g6777( .A1 (n6783), .A2 (y2079), .B (n6784), .Y (y3344) );
  OA21x2_ASAP7_75t_R   g6778( .A1 (n965), .A2 (n2163), .B (n2242), .Y (y3345) );
  AO21x1_ASAP7_75t_R   g6779( .A1 (n4273), .A2 (n22), .B (n529), .Y (n6787) );
  AO21x1_ASAP7_75t_R   g6780( .A1 (n5072), .A2 (n15), .B (n6787), .Y (y3346) );
  OA21x2_ASAP7_75t_R   g6781( .A1 (n103), .A2 (n116), .B (n123), .Y (y3347) );
  AND2x2_ASAP7_75t_R   g6782( .A (n466), .B (n604), .Y (y3348) );
  NOR2x1_ASAP7_75t_R   g6783( .A (n6443), .B (n6612), .Y (y3349) );
  AO21x1_ASAP7_75t_R   g6784( .A1 (n16), .A2 (n17), .B (n12), .Y (n6792) );
  NAND2x1_ASAP7_75t_R  g6785( .A (n6792), .B (n56), .Y (y3350) );
  OA21x2_ASAP7_75t_R   g6786( .A1 (n1537), .A2 (n1066), .B (n1641), .Y (y3351) );
  OA21x2_ASAP7_75t_R   g6787( .A1 (n1080), .A2 (n977), .B (n5942), .Y (y3353) );
  AO32x1_ASAP7_75t_R   g6788( .A1 (n3028), .A2 (n672), .A3 (n72), .B1 (y2079), .B2 (x4), .Y (y3354) );
  OR3x1_ASAP7_75t_R    g6789( .A (n529), .B (n3568), .C (n3294), .Y (y3355) );
  AO21x1_ASAP7_75t_R   g6790( .A1 (n360), .A2 (y2079), .B (x0), .Y (n6798) );
  OA21x2_ASAP7_75t_R   g6791( .A1 (n4250), .A2 (n12), .B (n6798), .Y (y3356) );
  AOI22x1_ASAP7_75t_R  g6792( .A1 (n22), .A2 (n3193), .B1 (x4), .B2 (n3004), .Y (y3357) );
  AND2x2_ASAP7_75t_R   g6793( .A (y1504), .B (n6643), .Y (y3358) );
  AND3x1_ASAP7_75t_R   g6794( .A (y2466), .B (n17), .C (x2), .Y (n6802) );
  INVx1_ASAP7_75t_R    g6795( .A (n6802), .Y (n6803) );
  AND2x2_ASAP7_75t_R   g6796( .A (n6803), .B (y1474), .Y (y3359) );
  AND2x2_ASAP7_75t_R   g6797( .A (n411), .B (n4619), .Y (y3360) );
  AND2x2_ASAP7_75t_R   g6798( .A (n3625), .B (y1474), .Y (y3361) );
  AND3x1_ASAP7_75t_R   g6799( .A (n3805), .B (n5910), .C (n4070), .Y (y3362) );
  NAND2x1_ASAP7_75t_R  g6800( .A (n17), .B (n4753), .Y (n6808) );
  INVx1_ASAP7_75t_R    g6801( .A (n6808), .Y (n6809) );
  AND2x2_ASAP7_75t_R   g6802( .A (y3758), .B (n1062), .Y (n6810) );
  AO21x1_ASAP7_75t_R   g6803( .A1 (n396), .A2 (n6809), .B (n6810), .Y (y3363) );
  AO21x1_ASAP7_75t_R   g6804( .A1 (y1757), .A2 (n125), .B (n4448), .Y (y3364) );
  OA21x2_ASAP7_75t_R   g6805( .A1 (n3005), .A2 (n22), .B (n5293), .Y (y3365) );
  NOR2x1_ASAP7_75t_R   g6806( .A (x2), .B (n1620), .Y (n6814) );
  INVx1_ASAP7_75t_R    g6807( .A (n6814), .Y (n6815) );
  OR3x1_ASAP7_75t_R    g6808( .A (y3758), .B (n5159), .C (n81), .Y (y3390) );
  AND2x2_ASAP7_75t_R   g6809( .A (n6815), .B (y3390), .Y (y3367) );
  AO21x1_ASAP7_75t_R   g6810( .A1 (n22), .A2 (n1572), .B (n3896), .Y (n6818) );
  AND3x1_ASAP7_75t_R   g6811( .A (n4876), .B (n3445), .C (y2079), .Y (n6819) );
  AO21x1_ASAP7_75t_R   g6812( .A1 (n4467), .A2 (n6818), .B (n6819), .Y (y3368) );
  INVx1_ASAP7_75t_R    g6813( .A (n4368), .Y (n6821) );
  AO21x1_ASAP7_75t_R   g6814( .A1 (n6821), .A2 (x5), .B (n5055), .Y (y3369) );
  AND2x2_ASAP7_75t_R   g6815( .A (n4441), .B (y3397), .Y (y3370) );
  AO21x1_ASAP7_75t_R   g6816( .A1 (n4632), .A2 (n4633), .B (n418), .Y (y3371) );
  AO21x1_ASAP7_75t_R   g6817( .A1 (n993), .A2 (n1469), .B (n2953), .Y (n6825) );
  AO21x1_ASAP7_75t_R   g6818( .A1 (n6825), .A2 (x0), .B (n2147), .Y (y3372) );
  AND2x2_ASAP7_75t_R   g6819( .A (n5059), .B (y3397), .Y (y3373) );
  OR3x1_ASAP7_75t_R    g6820( .A (n195), .B (n140), .C (n143), .Y (y3374) );
  OR3x1_ASAP7_75t_R    g6821( .A (n2964), .B (n6657), .C (n5323), .Y (y3375) );
  AND2x2_ASAP7_75t_R   g6822( .A (n4329), .B (y3397), .Y (y3376) );
  OR3x1_ASAP7_75t_R    g6823( .A (n1158), .B (n15), .C (n6306), .Y (n6831) );
  OR3x1_ASAP7_75t_R    g6824( .A (n3118), .B (y2466), .C (x2), .Y (n6832) );
  AND2x2_ASAP7_75t_R   g6825( .A (n6831), .B (n6832), .Y (y3378) );
  INVx1_ASAP7_75t_R    g6826( .A (n6698), .Y (n6834) );
  OA21x2_ASAP7_75t_R   g6827( .A1 (n3263), .A2 (n4108), .B (n6834), .Y (y3379) );
  AND2x2_ASAP7_75t_R   g6828( .A (n1064), .B (y648), .Y (y3380) );
  AND2x2_ASAP7_75t_R   g6829( .A (n1480), .B (x2), .Y (n6837) );
  XOR2x2_ASAP7_75t_R   g6830( .A (n2734), .B (n6837), .Y (y3381) );
  AO21x1_ASAP7_75t_R   g6831( .A1 (n22), .A2 (x5), .B (n211), .Y (n6839) );
  AO21x1_ASAP7_75t_R   g6832( .A1 (x4), .A2 (y2079), .B (n1838), .Y (n6840) );
  OA21x2_ASAP7_75t_R   g6833( .A1 (n4781), .A2 (n6839), .B (n6840), .Y (y3382) );
  AND2x2_ASAP7_75t_R   g6834( .A (y3397), .B (n3526), .Y (y3383) );
  OR3x1_ASAP7_75t_R    g6835( .A (n43), .B (n15), .C (n17), .Y (n6843) );
  AO21x1_ASAP7_75t_R   g6836( .A1 (n17), .A2 (n15), .B (n143), .Y (n6844) );
  INVx1_ASAP7_75t_R    g6837( .A (n6844), .Y (n6845) );
  OR3x1_ASAP7_75t_R    g6838( .A (n43), .B (x2), .C (x3), .Y (n6846) );
  INVx1_ASAP7_75t_R    g6839( .A (n6846), .Y (n6847) );
  AO21x1_ASAP7_75t_R   g6840( .A1 (n6843), .A2 (n6845), .B (n6847), .Y (n6848) );
  INVx1_ASAP7_75t_R    g6841( .A (n6848), .Y (y3384) );
  AND2x2_ASAP7_75t_R   g6842( .A (n411), .B (n3542), .Y (y3385) );
  OR3x1_ASAP7_75t_R    g6843( .A (n186), .B (y863), .C (n45), .Y (n6851) );
  AND2x2_ASAP7_75t_R   g6844( .A (n6747), .B (n6851), .Y (y3388) );
  AND2x2_ASAP7_75t_R   g6845( .A (n4545), .B (n3327), .Y (y3389) );
  AO21x1_ASAP7_75t_R   g6846( .A1 (n352), .A2 (n3085), .B (n3107), .Y (y3391) );
  AND2x2_ASAP7_75t_R   g6847( .A (n4651), .B (y3397), .Y (y3392) );
  INVx1_ASAP7_75t_R    g6848( .A (n948), .Y (n6856) );
  OR3x1_ASAP7_75t_R    g6849( .A (y3758), .B (n6856), .C (y863), .Y (y3393) );
  AO21x1_ASAP7_75t_R   g6850( .A1 (y9), .A2 (n418), .B (n1195), .Y (n6858) );
  XOR2x2_ASAP7_75t_R   g6851( .A (n6858), .B (x0), .Y (y3394) );
  AND3x1_ASAP7_75t_R   g6852( .A (n189), .B (n1319), .C (y2079), .Y (n6860) );
  AO21x1_ASAP7_75t_R   g6853( .A1 (n352), .A2 (n337), .B (n6860), .Y (y3395) );
  AND2x2_ASAP7_75t_R   g6854( .A (n4031), .B (n4633), .Y (y3396) );
  AND3x1_ASAP7_75t_R   g6855( .A (n315), .B (y2079), .C (n16), .Y (n6863) );
  NOR2x1_ASAP7_75t_R   g6856( .A (n392), .B (n6863), .Y (y3398) );
  AND3x1_ASAP7_75t_R   g6857( .A (y3293), .B (n3014), .C (x0), .Y (n6865) );
  INVx1_ASAP7_75t_R    g6858( .A (n6865), .Y (n6866) );
  AO21x1_ASAP7_75t_R   g6859( .A1 (n17), .A2 (x0), .B (n418), .Y (n6867) );
  AO21x1_ASAP7_75t_R   g6860( .A1 (x0), .A2 (y3293), .B (n6867), .Y (n6868) );
  AND2x2_ASAP7_75t_R   g6861( .A (n6866), .B (n6868), .Y (y3399) );
  AO21x1_ASAP7_75t_R   g6862( .A1 (n388), .A2 (n1163), .B (x3), .Y (n6870) );
  AO21x1_ASAP7_75t_R   g6863( .A1 (n310), .A2 (y2079), .B (n3338), .Y (n6871) );
  AND3x1_ASAP7_75t_R   g6864( .A (n6870), .B (n6871), .C (n1047), .Y (y3400) );
  AO21x1_ASAP7_75t_R   g6865( .A1 (y2079), .A2 (n22), .B (n45), .Y (n6873) );
  AO21x1_ASAP7_75t_R   g6866( .A1 (n1838), .A2 (y3293), .B (n6873), .Y (y3401) );
  AND3x1_ASAP7_75t_R   g6867( .A (n72), .B (n64), .C (n4976), .Y (y3402) );
  AND3x1_ASAP7_75t_R   g6868( .A (n3033), .B (n90), .C (n1295), .Y (n6876) );
  INVx1_ASAP7_75t_R    g6869( .A (n6876), .Y (n6877) );
  OA21x2_ASAP7_75t_R   g6870( .A1 (n2565), .A2 (n2545), .B (n6877), .Y (y3403) );
  NOR2x1_ASAP7_75t_R   g6871( .A (n392), .B (n4202), .Y (y3404) );
  AND2x2_ASAP7_75t_R   g6872( .A (y2578), .B (y1894), .Y (y3405) );
  AO21x1_ASAP7_75t_R   g6873( .A1 (n3040), .A2 (x5), .B (n347), .Y (n6881) );
  OA21x2_ASAP7_75t_R   g6874( .A1 (n4225), .A2 (n374), .B (y2079), .Y (n6882) );
  NOR2x1_ASAP7_75t_R   g6875( .A (n6881), .B (n6882), .Y (y3406) );
  AND2x2_ASAP7_75t_R   g6876( .A (n4107), .B (y2079), .Y (n6884) );
  OR3x1_ASAP7_75t_R    g6877( .A (n2964), .B (n6884), .C (n3263), .Y (y3407) );
  AND3x1_ASAP7_75t_R   g6878( .A (n380), .B (y1865), .C (n5819), .Y (y3408) );
  AO21x1_ASAP7_75t_R   g6879( .A1 (n5116), .A2 (x5), .B (n347), .Y (n6887) );
  INVx1_ASAP7_75t_R    g6880( .A (n6887), .Y (n6888) );
  AO21x1_ASAP7_75t_R   g6881( .A1 (n4129), .A2 (n6888), .B (n5998), .Y (y3409) );
  OR3x1_ASAP7_75t_R    g6882( .A (n347), .B (n12), .C (x5), .Y (n6890) );
  INVx1_ASAP7_75t_R    g6883( .A (n6890), .Y (n6891) );
  AO21x1_ASAP7_75t_R   g6884( .A1 (n382), .A2 (n685), .B (n6891), .Y (n6892) );
  AND2x2_ASAP7_75t_R   g6885( .A (n380), .B (n6892), .Y (y3410) );
  INVx1_ASAP7_75t_R    g6886( .A (n3457), .Y (n6894) );
  OA211x2_ASAP7_75t_R  g6887( .A1 (n6894), .A2 (n3502), .B (n1334), .C (y3852), .Y (y3411) );
  AND3x1_ASAP7_75t_R   g6888( .A (y3176), .B (n5493), .C (n652), .Y (y3412) );
  NAND2x1_ASAP7_75t_R  g6889( .A (n22), .B (n353), .Y (n6897) );
  OA21x2_ASAP7_75t_R   g6890( .A1 (n4360), .A2 (n22), .B (n6897), .Y (y3413) );
  AND2x2_ASAP7_75t_R   g6891( .A (y3172), .B (n3387), .Y (y3414) );
  AND2x2_ASAP7_75t_R   g6892( .A (n71), .B (n69), .Y (n6900) );
  AO21x1_ASAP7_75t_R   g6893( .A1 (n64), .A2 (n63), .B (n6900), .Y (y3415) );
  AND3x1_ASAP7_75t_R   g6894( .A (n84), .B (n125), .C (n22), .Y (n6902) );
  NAND2x1_ASAP7_75t_R  g6895( .A (y2079), .B (n6902), .Y (n6903) );
  AND2x2_ASAP7_75t_R   g6896( .A (n6903), .B (y1343), .Y (y3416) );
  AND3x1_ASAP7_75t_R   g6897( .A (n77), .B (n3804), .C (n4070), .Y (n6905) );
  INVx1_ASAP7_75t_R    g6898( .A (n6905), .Y (n6906) );
  OA21x2_ASAP7_75t_R   g6899( .A1 (x5), .A2 (n6906), .B (y2913), .Y (y3417) );
  OR3x1_ASAP7_75t_R    g6900( .A (y3758), .B (n4102), .C (n76), .Y (n6908) );
  NOR2x1_ASAP7_75t_R   g6901( .A (n17), .B (n3069), .Y (n6909) );
  INVx1_ASAP7_75t_R    g6902( .A (n6909), .Y (n6910) );
  NAND2x1_ASAP7_75t_R  g6903( .A (n6908), .B (n6910), .Y (y3418) );
  OR3x1_ASAP7_75t_R    g6904( .A (n145), .B (y2079), .C (x4), .Y (n6912) );
  OA21x2_ASAP7_75t_R   g6905( .A1 (n4360), .A2 (n22), .B (n6912), .Y (y3419) );
  NAND2x1_ASAP7_75t_R  g6906( .A (n4216), .B (n72), .Y (n6914) );
  INVx1_ASAP7_75t_R    g6907( .A (n6914), .Y (n6915) );
  AO21x1_ASAP7_75t_R   g6908( .A1 (n556), .A2 (n6915), .B (n4648), .Y (y3420) );
  AND2x2_ASAP7_75t_R   g6909( .A (n3647), .B (n685), .Y (y3421) );
  OR3x1_ASAP7_75t_R    g6910( .A (n987), .B (n143), .C (n529), .Y (y3422) );
  AO21x1_ASAP7_75t_R   g6911( .A1 (n559), .A2 (n310), .B (n1150), .Y (y3423) );
  OA21x2_ASAP7_75t_R   g6912( .A1 (n339), .A2 (n403), .B (n3119), .Y (y3424) );
  AND3x1_ASAP7_75t_R   g6913( .A (n413), .B (n724), .C (y3377), .Y (y3425) );
  AO21x1_ASAP7_75t_R   g6914( .A1 (n6821), .A2 (x5), .B (n2051), .Y (y3426) );
  AO32x1_ASAP7_75t_R   g6915( .A1 (y1281), .A2 (n451), .A3 (x3), .B1 (x5), .B2 (n2994), .Y (y3429) );
  AO32x1_ASAP7_75t_R   g6916( .A1 (y3852), .A2 (n90), .A3 (n1502), .B1 (n15), .B2 (n1245), .Y (y3430) );
  OA21x2_ASAP7_75t_R   g6917( .A1 (n4920), .A2 (n3376), .B (n4507), .Y (y3431) );
  NAND2x1_ASAP7_75t_R  g6918( .A (y2079), .B (n910), .Y (n6926) );
  INVx1_ASAP7_75t_R    g6919( .A (n6926), .Y (y3432) );
  AND3x1_ASAP7_75t_R   g6920( .A (n537), .B (n17), .C (x5), .Y (n6928) );
  AO21x1_ASAP7_75t_R   g6921( .A1 (n5373), .A2 (n556), .B (n6928), .Y (y3433) );
  AO21x1_ASAP7_75t_R   g6922( .A1 (y19), .A2 (n52), .B (n53), .Y (y3434) );
  AND2x2_ASAP7_75t_R   g6923( .A (n113), .B (x3), .Y (n6931) );
  AO21x1_ASAP7_75t_R   g6924( .A1 (n17), .A2 (n747), .B (n6931), .Y (y3435) );
  NAND2x1_ASAP7_75t_R  g6925( .A (x5), .B (n974), .Y (n6933) );
  INVx1_ASAP7_75t_R    g6926( .A (n6933), .Y (n6934) );
  AO21x1_ASAP7_75t_R   g6927( .A1 (n1196), .A2 (y1894), .B (n6934), .Y (y3436) );
  AND3x1_ASAP7_75t_R   g6928( .A (n4116), .B (n310), .C (n388), .Y (n6936) );
  AO21x1_ASAP7_75t_R   g6929( .A1 (n556), .A2 (n5373), .B (n6936), .Y (y3437) );
  OR3x1_ASAP7_75t_R    g6930( .A (n581), .B (n1137), .C (n344), .Y (y3438) );
  NAND2x1_ASAP7_75t_R  g6931( .A (n4526), .B (n2992), .Y (y3439) );
  OA21x2_ASAP7_75t_R   g6932( .A1 (x3), .A2 (n1927), .B (n5843), .Y (y3440) );
  AO21x1_ASAP7_75t_R   g6933( .A1 (n388), .A2 (n310), .B (x3), .Y (n6941) );
  AND2x2_ASAP7_75t_R   g6934( .A (n5843), .B (n6941), .Y (y3441) );
  AND3x1_ASAP7_75t_R   g6935( .A (n3109), .B (y3176), .C (n348), .Y (y3442) );
  INVx1_ASAP7_75t_R    g6936( .A (n6881), .Y (n6944) );
  OA21x2_ASAP7_75t_R   g6937( .A1 (y2347), .A2 (n6944), .B (n380), .Y (y3443) );
  AND2x2_ASAP7_75t_R   g6938( .A (n5843), .B (n3648), .Y (y3444) );
  OA21x2_ASAP7_75t_R   g6939( .A1 (n503), .A2 (n1948), .B (n219), .Y (y3446) );
  AO21x1_ASAP7_75t_R   g6940( .A1 (n3269), .A2 (n660), .B (n3443), .Y (y3448) );
  AND2x2_ASAP7_75t_R   g6941( .A (y2424), .B (n348), .Y (y3449) );
  OR3x1_ASAP7_75t_R    g6942( .A (n628), .B (n2994), .C (n3080), .Y (y3450) );
  AO21x1_ASAP7_75t_R   g6943( .A1 (n1047), .A2 (n1082), .B (n1075), .Y (y3451) );
  INVx1_ASAP7_75t_R    g6944( .A (n191), .Y (n6952) );
  AO21x1_ASAP7_75t_R   g6945( .A1 (n6952), .A2 (n16), .B (n2169), .Y (n6953) );
  XOR2x2_ASAP7_75t_R   g6946( .A (n6953), .B (n17), .Y (y3452) );
  AO32x1_ASAP7_75t_R   g6947( .A1 (n22), .A2 (n316), .A3 (n397), .B1 (x4), .B2 (n3193), .Y (y3453) );
  AND2x2_ASAP7_75t_R   g6948( .A (y3176), .B (n5493), .Y (y3454) );
  AND2x2_ASAP7_75t_R   g6949( .A (n3256), .B (n5843), .Y (y3455) );
  NAND2x1_ASAP7_75t_R  g6950( .A (x4), .B (n2997), .Y (n6958) );
  AND2x2_ASAP7_75t_R   g6951( .A (n3987), .B (n6958), .Y (y3456) );
  NOR2x1_ASAP7_75t_R   g6952( .A (n15), .B (n143), .Y (n6960) );
  NOR2x1_ASAP7_75t_R   g6953( .A (n2164), .B (n6960), .Y (y3457) );
  NOR2x1_ASAP7_75t_R   g6954( .A (n3747), .B (n1927), .Y (y3458) );
  AO21x1_ASAP7_75t_R   g6955( .A1 (n342), .A2 (n17), .B (n293), .Y (y3459) );
  INVx1_ASAP7_75t_R    g6956( .A (y2584), .Y (n6964) );
  AND3x1_ASAP7_75t_R   g6957( .A (n6964), .B (y193), .C (y3808), .Y (y3460) );
  NAND2x1_ASAP7_75t_R  g6958( .A (x5), .B (n3978), .Y (n6966) );
  AND2x2_ASAP7_75t_R   g6959( .A (n6173), .B (n6966), .Y (y3461) );
  OA211x2_ASAP7_75t_R  g6960( .A1 (n718), .A2 (n4116), .B (n3326), .C (n84), .Y (y3462) );
  INVx1_ASAP7_75t_R    g6961( .A (n1587), .Y (y3463) );
  OR3x1_ASAP7_75t_R    g6962( .A (n418), .B (n12), .C (x3), .Y (n6970) );
  INVx1_ASAP7_75t_R    g6963( .A (n6970), .Y (n6971) );
  AO21x1_ASAP7_75t_R   g6964( .A1 (n28), .A2 (n388), .B (n125), .Y (n6972) );
  OA21x2_ASAP7_75t_R   g6965( .A1 (y2626), .A2 (n6971), .B (n6972), .Y (y3464) );
  AND3x1_ASAP7_75t_R   g6966( .A (n4039), .B (n4619), .C (n4618), .Y (y3465) );
  AND2x2_ASAP7_75t_R   g6967( .A (n3426), .B (n84), .Y (n6975) );
  AO21x1_ASAP7_75t_R   g6968( .A1 (n6975), .A2 (n6609), .B (n6928), .Y (y3466) );
  AO21x1_ASAP7_75t_R   g6969( .A1 (n310), .A2 (x3), .B (n3386), .Y (n6977) );
  NOR2x1_ASAP7_75t_R   g6970( .A (y2079), .B (n2992), .Y (n6978) );
  AO21x1_ASAP7_75t_R   g6971( .A1 (y2079), .A2 (n6977), .B (n6978), .Y (y3467) );
  AND3x1_ASAP7_75t_R   g6972( .A (n3326), .B (n6466), .C (n387), .Y (y3468) );
  AO21x1_ASAP7_75t_R   g6973( .A1 (n12), .A2 (n20), .B (y269), .Y (y3469) );
  AO21x1_ASAP7_75t_R   g6974( .A1 (n16), .A2 (n1186), .B (n1083), .Y (y3470) );
  NOR2x1_ASAP7_75t_R   g6975( .A (n12), .B (n3118), .Y (n6983) );
  OA21x2_ASAP7_75t_R   g6976( .A1 (n337), .A2 (n6983), .B (n4016), .Y (y3471) );
  NAND2x1_ASAP7_75t_R  g6977( .A (n5256), .B (n28), .Y (n6985) );
  AO32x1_ASAP7_75t_R   g6978( .A1 (n28), .A2 (n5256), .A3 (n6230), .B1 (n6985), .B2 (n6229), .Y (y3472) );
  AO21x1_ASAP7_75t_R   g6979( .A1 (y1693), .A2 (x0), .B (n630), .Y (y3473) );
  INVx1_ASAP7_75t_R    g6980( .A (n1175), .Y (n6988) );
  INVx1_ASAP7_75t_R    g6981( .A (n690), .Y (n6989) );
  AO221x2_ASAP7_75t_R  g6982( .A1 (n6988), .A2 (n6989), .B1 (n1175), .B2 (n690), .C (n143), .Y (y3474) );
  AND3x1_ASAP7_75t_R   g6983( .A (n369), .B (n388), .C (n12), .Y (n6991) );
  NOR2x1_ASAP7_75t_R   g6984( .A (n3118), .B (n6991), .Y (y3475) );
  AND3x1_ASAP7_75t_R   g6985( .A (n3882), .B (n3387), .C (n299), .Y (y3476) );
  AO21x1_ASAP7_75t_R   g6986( .A1 (y2079), .A2 (x3), .B (n315), .Y (n6994) );
  AO21x1_ASAP7_75t_R   g6987( .A1 (n360), .A2 (n6994), .B (n5631), .Y (y3477) );
  OR3x1_ASAP7_75t_R    g6988( .A (n2001), .B (n3417), .C (n143), .Y (y3478) );
  AO32x1_ASAP7_75t_R   g6989( .A1 (n22), .A2 (n397), .A3 (n4451), .B1 (x4), .B2 (n3193), .Y (y3479) );
  AO21x1_ASAP7_75t_R   g6990( .A1 (n527), .A2 (n765), .B (n957), .Y (y3480) );
  AND2x2_ASAP7_75t_R   g6991( .A (n330), .B (x5), .Y (n6999) );
  OA21x2_ASAP7_75t_R   g6992( .A1 (n377), .A2 (n6999), .B (n5727), .Y (y3481) );
  INVx1_ASAP7_75t_R    g6993( .A (n5507), .Y (n7001) );
  NOR2x1_ASAP7_75t_R   g6994( .A (n7001), .B (n4768), .Y (y3482) );
  AO21x1_ASAP7_75t_R   g6995( .A1 (n3023), .A2 (n3776), .B (n3279), .Y (y3483) );
  AND2x2_ASAP7_75t_R   g6996( .A (y2701), .B (n5479), .Y (y3484) );
  AO21x1_ASAP7_75t_R   g6997( .A1 (n310), .A2 (y2068), .B (n6978), .Y (y3485) );
  AO21x1_ASAP7_75t_R   g6998( .A1 (n3354), .A2 (y3293), .B (x0), .Y (y3486) );
  OA21x2_ASAP7_75t_R   g6999( .A1 (n3193), .A2 (n3085), .B (n5342), .Y (y3487) );
  OA211x2_ASAP7_75t_R  g7000( .A1 (n408), .A2 (n529), .B (n6941), .C (n3884), .Y (y3488) );
  AO21x1_ASAP7_75t_R   g7001( .A1 (n455), .A2 (n45), .B (n3298), .Y (y3489) );
  AO21x1_ASAP7_75t_R   g7002( .A1 (n481), .A2 (n660), .B (y2196), .Y (n7010) );
  XOR2x2_ASAP7_75t_R   g7003( .A (n7010), .B (n378), .Y (y3490) );
  AO21x1_ASAP7_75t_R   g7004( .A1 (y1281), .A2 (x3), .B (n6367), .Y (y3491) );
  AND2x2_ASAP7_75t_R   g7005( .A (n397), .B (n22), .Y (n7013) );
  OA21x2_ASAP7_75t_R   g7006( .A1 (n3193), .A2 (n7013), .B (n4835), .Y (y3492) );
  NOR2x1_ASAP7_75t_R   g7007( .A (n300), .B (n4282), .Y (n7015) );
  OA21x2_ASAP7_75t_R   g7008( .A1 (n7015), .A2 (x3), .B (n3882), .Y (y3493) );
  AND3x1_ASAP7_75t_R   g7009( .A (n776), .B (n388), .C (n12), .Y (n7017) );
  AO21x1_ASAP7_75t_R   g7010( .A1 (n25), .A2 (x0), .B (n7017), .Y (y3494) );
  INVx1_ASAP7_75t_R    g7011( .A (n5513), .Y (n7019) );
  AO21x1_ASAP7_75t_R   g7012( .A1 (n7019), .A2 (n299), .B (y2079), .Y (y3514) );
  AND2x2_ASAP7_75t_R   g7013( .A (n5514), .B (y3514), .Y (y3495) );
  AND2x2_ASAP7_75t_R   g7014( .A (y271), .B (n1310), .Y (y3496) );
  AND2x2_ASAP7_75t_R   g7015( .A (n6344), .B (n3648), .Y (y3497) );
  OA21x2_ASAP7_75t_R   g7016( .A1 (n4584), .A2 (y1300), .B (n3648), .Y (y3498) );
  INVx1_ASAP7_75t_R    g7017( .A (n1166), .Y (n7025) );
  INVx1_ASAP7_75t_R    g7018( .A (n1186), .Y (n7026) );
  AO21x1_ASAP7_75t_R   g7019( .A1 (n7026), .A2 (n1166), .B (n529), .Y (y3980) );
  AO21x1_ASAP7_75t_R   g7020( .A1 (n7025), .A2 (n1186), .B (y3980), .Y (y3499) );
  AO21x1_ASAP7_75t_R   g7021( .A1 (n2246), .A2 (n4336), .B (n6928), .Y (y3500) );
  AO21x1_ASAP7_75t_R   g7022( .A1 (y2079), .A2 (n3325), .B (n914), .Y (n7030) );
  AO21x1_ASAP7_75t_R   g7023( .A1 (n7030), .A2 (n4583), .B (n6367), .Y (y3501) );
  AO21x1_ASAP7_75t_R   g7024( .A1 (n111), .A2 (n15), .B (n146), .Y (y3502) );
  NAND2x1_ASAP7_75t_R  g7025( .A (n1536), .B (n2848), .Y (n7033) );
  AND2x2_ASAP7_75t_R   g7026( .A (n7033), .B (n4261), .Y (y3503) );
  OA33x2_ASAP7_75t_R   g7027( .A1 (x4), .A2 (n303), .A3 (n145), .B1 (n628), .B2 (n22), .B3 (n2718), .Y (y3504) );
  AND2x2_ASAP7_75t_R   g7028( .A (n4016), .B (n922), .Y (y3505) );
  INVx1_ASAP7_75t_R    g7029( .A (n897), .Y (n7037) );
  AND2x2_ASAP7_75t_R   g7030( .A (n2825), .B (n52), .Y (n7038) );
  AND3x1_ASAP7_75t_R   g7031( .A (n1676), .B (n17), .C (x0), .Y (n7039) );
  INVx1_ASAP7_75t_R    g7032( .A (n7039), .Y (n7040) );
  OA21x2_ASAP7_75t_R   g7033( .A1 (n7037), .A2 (n7038), .B (n7040), .Y (y3506) );
  NOR2x1_ASAP7_75t_R   g7034( .A (n368), .B (n3370), .Y (n7042) );
  AO21x1_ASAP7_75t_R   g7035( .A1 (n125), .A2 (n3085), .B (n7042), .Y (y3507) );
  INVx1_ASAP7_75t_R    g7036( .A (n2848), .Y (n7044) );
  OA21x2_ASAP7_75t_R   g7037( .A1 (n7044), .A2 (n2315), .B (n2729), .Y (y3508) );
  AO21x1_ASAP7_75t_R   g7038( .A1 (n137), .A2 (n72), .B (n518), .Y (n7046) );
  OA21x2_ASAP7_75t_R   g7039( .A1 (n218), .A2 (n3446), .B (n7046), .Y (y3509) );
  AO21x1_ASAP7_75t_R   g7040( .A1 (n12), .A2 (n17), .B (y2079), .Y (n7048) );
  AO21x1_ASAP7_75t_R   g7041( .A1 (n377), .A2 (n7048), .B (n6821), .Y (y3510) );
  AND2x2_ASAP7_75t_R   g7042( .A (n2984), .B (n3882), .Y (y3511) );
  AND2x2_ASAP7_75t_R   g7043( .A (n4016), .B (y2727), .Y (y3512) );
  AND2x2_ASAP7_75t_R   g7044( .A (y2727), .B (n3387), .Y (y3513) );
  AND3x1_ASAP7_75t_R   g7045( .A (n323), .B (n388), .C (n360), .Y (n7053) );
  INVx1_ASAP7_75t_R    g7046( .A (n7053), .Y (n7054) );
  NOR2x1_ASAP7_75t_R   g7047( .A (x5), .B (x3), .Y (n7055) );
  AO21x1_ASAP7_75t_R   g7048( .A1 (n7055), .A2 (n22), .B (x0), .Y (n7056) );
  AND2x2_ASAP7_75t_R   g7049( .A (n7054), .B (n7056), .Y (y3515) );
  AND2x2_ASAP7_75t_R   g7050( .A (n3600), .B (y1894), .Y (y3516) );
  AND2x2_ASAP7_75t_R   g7051( .A (y3172), .B (n3797), .Y (y3517) );
  AO21x1_ASAP7_75t_R   g7052( .A1 (n1158), .A2 (y2079), .B (x0), .Y (n7060) );
  AND2x2_ASAP7_75t_R   g7053( .A (n7060), .B (n4618), .Y (y3518) );
  AO21x1_ASAP7_75t_R   g7054( .A1 (n740), .A2 (n337), .B (n628), .Y (y3519) );
  NOR2x1_ASAP7_75t_R   g7055( .A (n1160), .B (n481), .Y (n7063) );
  AND2x2_ASAP7_75t_R   g7056( .A (n3647), .B (n7063), .Y (y3520) );
  OAI21x1_ASAP7_75t_R  g7057( .A1 (n6134), .A2 (n12), .B (y2516), .Y (y3521) );
  AO21x1_ASAP7_75t_R   g7058( .A1 (n5520), .A2 (n1572), .B (y2079), .Y (y3522) );
  NAND2x1_ASAP7_75t_R  g7059( .A (n12), .B (n285), .Y (n7067) );
  AND2x2_ASAP7_75t_R   g7060( .A (n3647), .B (n7067), .Y (y3523) );
  AND2x2_ASAP7_75t_R   g7061( .A (y2727), .B (n645), .Y (y3524) );
  AO21x1_ASAP7_75t_R   g7062( .A1 (n1572), .A2 (n5520), .B (n529), .Y (y3525) );
  AO21x1_ASAP7_75t_R   g7063( .A1 (n4225), .A2 (x5), .B (n349), .Y (y3526) );
  AO21x1_ASAP7_75t_R   g7064( .A1 (x5), .A2 (n4225), .B (n2051), .Y (y3528) );
  AO21x1_ASAP7_75t_R   g7065( .A1 (n178), .A2 (n67), .B (n13), .Y (y3529) );
  NOR2x1_ASAP7_75t_R   g7066( .A (n756), .B (n3360), .Y (n7074) );
  NOR2x1_ASAP7_75t_R   g7067( .A (n4340), .B (n7074), .Y (y3530) );
  AO21x1_ASAP7_75t_R   g7068( .A1 (x5), .A2 (n3414), .B (n676), .Y (y3531) );
  OA21x2_ASAP7_75t_R   g7069( .A1 (n2994), .A2 (n3426), .B (n3391), .Y (y3532) );
  AO21x1_ASAP7_75t_R   g7070( .A1 (n1903), .A2 (y3852), .B (n990), .Y (y3533) );
  OR3x1_ASAP7_75t_R    g7071( .A (y772), .B (n2001), .C (n1907), .Y (y3534) );
  AND3x1_ASAP7_75t_R   g7072( .A (n5843), .B (n451), .C (n4508), .Y (y3535) );
  AND2x2_ASAP7_75t_R   g7073( .A (y1693), .B (n1342), .Y (y3536) );
  AO21x1_ASAP7_75t_R   g7074( .A1 (n3284), .A2 (x0), .B (n3443), .Y (y3537) );
  AND2x2_ASAP7_75t_R   g7075( .A (n5843), .B (n4508), .Y (y3538) );
  AO21x1_ASAP7_75t_R   g7076( .A1 (x1), .A2 (n2590), .B (n2546), .Y (y3539) );
  INVx1_ASAP7_75t_R    g7077( .A (n5641), .Y (n7085) );
  AO21x1_ASAP7_75t_R   g7078( .A1 (n348), .A2 (n5055), .B (n7085), .Y (y3540) );
  AND2x2_ASAP7_75t_R   g7079( .A (n2282), .B (n1490), .Y (y3541) );
  AND3x1_ASAP7_75t_R   g7080( .A (y1903), .B (n645), .C (n1851), .Y (y3542) );
  AO21x1_ASAP7_75t_R   g7081( .A1 (y2079), .A2 (n3384), .B (n5403), .Y (y3543) );
  OR3x1_ASAP7_75t_R    g7082( .A (n2995), .B (n6928), .C (n3574), .Y (y3544) );
  AND2x2_ASAP7_75t_R   g7083( .A (n3497), .B (n556), .Y (y3545) );
  AO21x1_ASAP7_75t_R   g7084( .A1 (y2079), .A2 (n3792), .B (n5403), .Y (y3546) );
  AND2x2_ASAP7_75t_R   g7085( .A (n5843), .B (n645), .Y (y3547) );
  AO21x1_ASAP7_75t_R   g7086( .A1 (y2079), .A2 (n3325), .B (n5403), .Y (y3548) );
  AND2x2_ASAP7_75t_R   g7087( .A (y2754), .B (n1334), .Y (y3549) );
  AO21x1_ASAP7_75t_R   g7088( .A1 (n495), .A2 (x2), .B (x0), .Y (y3550) );
  OA21x2_ASAP7_75t_R   g7089( .A1 (n4702), .A2 (y772), .B (n2701), .Y (y3551) );
  AO21x1_ASAP7_75t_R   g7090( .A1 (n3284), .A2 (x0), .B (n4541), .Y (y3552) );
  INVx1_ASAP7_75t_R    g7091( .A (n3436), .Y (n7099) );
  AND3x1_ASAP7_75t_R   g7092( .A (n7099), .B (n84), .C (n556), .Y (y3553) );
  AND2x2_ASAP7_75t_R   g7093( .A (n6159), .B (n1342), .Y (y3554) );
  AND3x1_ASAP7_75t_R   g7094( .A (n6033), .B (n3943), .C (n556), .Y (y3555) );
  NOR2x1_ASAP7_75t_R   g7095( .A (n65), .B (n1514), .Y (y3557) );
  AO21x1_ASAP7_75t_R   g7096( .A1 (n6190), .A2 (x0), .B (n628), .Y (y3558) );
  NOR2x1_ASAP7_75t_R   g7097( .A (n5994), .B (n4486), .Y (y3559) );
  AO21x1_ASAP7_75t_R   g7098( .A1 (n6190), .A2 (x0), .B (n3415), .Y (y3560) );
  AND3x1_ASAP7_75t_R   g7099( .A (n3027), .B (x5), .C (x3), .Y (n7107) );
  INVx1_ASAP7_75t_R    g7100( .A (n7107), .Y (n7108) );
  OR3x1_ASAP7_75t_R    g7101( .A (n211), .B (x4), .C (x5), .Y (n7109) );
  AND3x1_ASAP7_75t_R   g7102( .A (n7108), .B (n7109), .C (n1062), .Y (y3561) );
  AND2x2_ASAP7_75t_R   g7103( .A (n2182), .B (n2701), .Y (y3562) );
  NAND2x1_ASAP7_75t_R  g7104( .A (n334), .B (n4526), .Y (y3563) );
  AO21x1_ASAP7_75t_R   g7105( .A1 (x5), .A2 (n4225), .B (n286), .Y (y3564) );
  NOR2x1_ASAP7_75t_R   g7106( .A (n12), .B (y2466), .Y (n7114) );
  AO21x1_ASAP7_75t_R   g7107( .A1 (n382), .A2 (n7114), .B (n6253), .Y (y3565) );
  OR3x1_ASAP7_75t_R    g7108( .A (y1081), .B (n787), .C (n109), .Y (y3566) );
  NAND2x1_ASAP7_75t_R  g7109( .A (n12), .B (n883), .Y (n7117) );
  AO21x1_ASAP7_75t_R   g7110( .A1 (n806), .A2 (n7117), .B (n81), .Y (y3567) );
  OA21x2_ASAP7_75t_R   g7111( .A1 (n2534), .A2 (n276), .B (n64), .Y (y3568) );
  OA21x2_ASAP7_75t_R   g7112( .A1 (n231), .A2 (n1851), .B (n3176), .Y (y3569) );
  OA21x2_ASAP7_75t_R   g7113( .A1 (n421), .A2 (n1851), .B (n556), .Y (y3570) );
  AO21x1_ASAP7_75t_R   g7114( .A1 (n413), .A2 (n348), .B (x5), .Y (n7122) );
  AND2x2_ASAP7_75t_R   g7115( .A (n7122), .B (y2727), .Y (y3571) );
  AND2x2_ASAP7_75t_R   g7116( .A (y168), .B (n672), .Y (y3572) );
  AO21x1_ASAP7_75t_R   g7117( .A1 (y2079), .A2 (n22), .B (y2998), .Y (y3573) );
  NAND2x1_ASAP7_75t_R  g7118( .A (n4708), .B (n5127), .Y (n7126) );
  OA21x2_ASAP7_75t_R   g7119( .A1 (n4317), .A2 (x5), .B (n7126), .Y (y3574) );
  AO21x1_ASAP7_75t_R   g7120( .A1 (n765), .A2 (n1952), .B (n1140), .Y (y3575) );
  AO21x1_ASAP7_75t_R   g7121( .A1 (y2079), .A2 (x0), .B (n403), .Y (n7129) );
  INVx1_ASAP7_75t_R    g7122( .A (n7129), .Y (n7130) );
  INVx1_ASAP7_75t_R    g7123( .A (n6019), .Y (n7131) );
  AO21x1_ASAP7_75t_R   g7124( .A1 (y168), .A2 (n7130), .B (n7131), .Y (y3576) );
  OR3x1_ASAP7_75t_R    g7125( .A (n1032), .B (x4), .C (x5), .Y (n7133) );
  AND2x2_ASAP7_75t_R   g7126( .A (n7133), .B (n4959), .Y (n7134) );
  NAND2x1_ASAP7_75t_R  g7127( .A (x5), .B (n409), .Y (n7135) );
  OA21x2_ASAP7_75t_R   g7128( .A1 (n7134), .A2 (x0), .B (n7135), .Y (y3577) );
  AND2x2_ASAP7_75t_R   g7129( .A (n67), .B (y2079), .Y (n7137) );
  AO21x1_ASAP7_75t_R   g7130( .A1 (x1), .A2 (n2210), .B (n7137), .Y (y3578) );
  AND2x2_ASAP7_75t_R   g7131( .A (y1903), .B (n3139), .Y (y3579) );
  AND2x2_ASAP7_75t_R   g7132( .A (n1881), .B (n968), .Y (y3580) );
  OA21x2_ASAP7_75t_R   g7133( .A1 (n2164), .A2 (x0), .B (n2836), .Y (y3581) );
  AND2x2_ASAP7_75t_R   g7134( .A (n4171), .B (y2319), .Y (y3582) );
  OA21x2_ASAP7_75t_R   g7135( .A1 (n3039), .A2 (n58), .B (n5828), .Y (y3583) );
  AO21x1_ASAP7_75t_R   g7136( .A1 (y2079), .A2 (n948), .B (n2107), .Y (n7144) );
  AND3x1_ASAP7_75t_R   g7137( .A (n231), .B (n22), .C (n12), .Y (n7145) );
  INVx1_ASAP7_75t_R    g7138( .A (n7145), .Y (n7146) );
  OA21x2_ASAP7_75t_R   g7139( .A1 (n7144), .A2 (y863), .B (n7146), .Y (y3584) );
  AND3x1_ASAP7_75t_R   g7140( .A (n299), .B (n408), .C (x5), .Y (n7148) );
  AO21x1_ASAP7_75t_R   g7141( .A1 (x3), .A2 (n1775), .B (n7148), .Y (y3585) );
  AO21x1_ASAP7_75t_R   g7142( .A1 (n310), .A2 (y2068), .B (n6690), .Y (y3586) );
  AO32x1_ASAP7_75t_R   g7143( .A1 (n17), .A2 (n352), .A3 (n3480), .B1 (n3457), .B2 (y104), .Y (y3587) );
  NAND2x1_ASAP7_75t_R  g7144( .A (y3377), .B (n686), .Y (n7152) );
  AND2x2_ASAP7_75t_R   g7145( .A (n7152), .B (n5828), .Y (y3588) );
  AO21x1_ASAP7_75t_R   g7146( .A1 (n2825), .A2 (n52), .B (n1317), .Y (y3589) );
  AO21x1_ASAP7_75t_R   g7147( .A1 (n16), .A2 (x5), .B (y2022), .Y (n7155) );
  AO21x1_ASAP7_75t_R   g7148( .A1 (n7155), .A2 (n15), .B (n2156), .Y (y3590) );
  OA21x2_ASAP7_75t_R   g7149( .A1 (n6977), .A2 (n7026), .B (n3882), .Y (y3591) );
  AO32x1_ASAP7_75t_R   g7150( .A1 (n556), .A2 (n125), .A3 (n3457), .B1 (x5), .B2 (n3521), .Y (y3592) );
  NOR2x1_ASAP7_75t_R   g7151( .A (n518), .B (n5372), .Y (n7159) );
  OR3x1_ASAP7_75t_R    g7152( .A (n7159), .B (n3192), .C (n630), .Y (y3593) );
  AO21x1_ASAP7_75t_R   g7153( .A1 (y2079), .A2 (x0), .B (n4514), .Y (y3594) );
  AO21x1_ASAP7_75t_R   g7154( .A1 (n22), .A2 (x0), .B (n3443), .Y (n7162) );
  AO21x1_ASAP7_75t_R   g7155( .A1 (n421), .A2 (n299), .B (n7162), .Y (y3595) );
  AO32x1_ASAP7_75t_R   g7156( .A1 (n388), .A2 (n84), .A3 (n3128), .B1 (x4), .B2 (n628), .Y (y3596) );
  OR3x1_ASAP7_75t_R    g7157( .A (n6690), .B (n628), .C (n630), .Y (y3597) );
  AO21x1_ASAP7_75t_R   g7158( .A1 (n3109), .A2 (y3176), .B (n347), .Y (y3599) );
  NAND2x1_ASAP7_75t_R  g7159( .A (n473), .B (n299), .Y (n7167) );
  AND2x2_ASAP7_75t_R   g7160( .A (n7167), .B (n17), .Y (n7168) );
  NOR2x1_ASAP7_75t_R   g7161( .A (n5894), .B (n7168), .Y (y3600) );
  AO21x1_ASAP7_75t_R   g7162( .A1 (y1300), .A2 (n3325), .B (n4584), .Y (y3601) );
  AND2x2_ASAP7_75t_R   g7163( .A (n67), .B (n1510), .Y (y3603) );
  AO21x1_ASAP7_75t_R   g7164( .A1 (n3013), .A2 (n419), .B (n17), .Y (n7172) );
  AND2x2_ASAP7_75t_R   g7165( .A (n7172), .B (n1062), .Y (y3604) );
  AO21x1_ASAP7_75t_R   g7166( .A1 (n3469), .A2 (n5385), .B (n3472), .Y (y3605) );
  AND2x2_ASAP7_75t_R   g7167( .A (y1903), .B (n401), .Y (y3606) );
  AO21x1_ASAP7_75t_R   g7168( .A1 (n2246), .A2 (n4336), .B (n3192), .Y (y3607) );
  NAND2x1_ASAP7_75t_R  g7169( .A (n334), .B (n316), .Y (y3608) );
  AO32x1_ASAP7_75t_R   g7170( .A1 (x3), .A2 (n3013), .A3 (n419), .B1 (n17), .B2 (n3823), .Y (y3609) );
  AO21x1_ASAP7_75t_R   g7171( .A1 (n72), .A2 (n64), .B (n145), .Y (y3610) );
  AND2x2_ASAP7_75t_R   g7172( .A (n4111), .B (y2727), .Y (y3611) );
  AO32x1_ASAP7_75t_R   g7173( .A1 (x5), .A2 (n72), .A3 (n4551), .B1 (y2079), .B2 (n3629), .Y (y3612) );
  NAND2x1_ASAP7_75t_R  g7174( .A (x5), .B (n3325), .Y (n7182) );
  AO21x1_ASAP7_75t_R   g7175( .A1 (n4111), .A2 (n7182), .B (n914), .Y (y3613) );
  AND3x1_ASAP7_75t_R   g7176( .A (n3477), .B (n5828), .C (n724), .Y (y3614) );
  NOR2x1_ASAP7_75t_R   g7177( .A (n17), .B (n3027), .Y (n7185) );
  AO21x1_ASAP7_75t_R   g7178( .A1 (n369), .A2 (x2), .B (n7185), .Y (y3615) );
  AO21x1_ASAP7_75t_R   g7179( .A1 (n645), .A2 (n3085), .B (n7042), .Y (y3616) );
  INVx1_ASAP7_75t_R    g7180( .A (n1466), .Y (n7188) );
  AO21x1_ASAP7_75t_R   g7181( .A1 (n1337), .A2 (n7188), .B (y773), .Y (y3617) );
  AO21x1_ASAP7_75t_R   g7182( .A1 (n72), .A2 (n529), .B (n4420), .Y (y3618) );
  AO21x1_ASAP7_75t_R   g7183( .A1 (n382), .A2 (x0), .B (y2723), .Y (y3619) );
  OR3x1_ASAP7_75t_R    g7184( .A (n3095), .B (n2994), .C (n628), .Y (y3620) );
  OA21x2_ASAP7_75t_R   g7185( .A1 (x3), .A2 (n1137), .B (n4755), .Y (y3621) );
  AO21x1_ASAP7_75t_R   g7186( .A1 (n1255), .A2 (x2), .B (n61), .Y (n7194) );
  XOR2x2_ASAP7_75t_R   g7187( .A (n7194), .B (n17), .Y (y3622) );
  INVx1_ASAP7_75t_R    g7188( .A (n3325), .Y (n7196) );
  AND3x1_ASAP7_75t_R   g7189( .A (n7196), .B (n352), .C (n28), .Y (n7197) );
  INVx1_ASAP7_75t_R    g7190( .A (n7197), .Y (n7198) );
  NAND2x1_ASAP7_75t_R  g7191( .A (n5800), .B (n7198), .Y (y3623) );
  AO21x1_ASAP7_75t_R   g7192( .A1 (n16), .A2 (n2514), .B (n2527), .Y (y3624) );
  OA21x2_ASAP7_75t_R   g7193( .A1 (n5678), .A2 (n4052), .B (n4633), .Y (y3625) );
  NAND2x1_ASAP7_75t_R  g7194( .A (n22), .B (n3645), .Y (n7202) );
  AND3x1_ASAP7_75t_R   g7195( .A (y1903), .B (n7202), .C (n672), .Y (y3626) );
  AO21x1_ASAP7_75t_R   g7196( .A1 (n178), .A2 (x0), .B (n182), .Y (y3627) );
  OR3x1_ASAP7_75t_R    g7197( .A (n315), .B (n403), .C (x5), .Y (n7205) );
  OA21x2_ASAP7_75t_R   g7198( .A1 (n6610), .A2 (y2079), .B (n7205), .Y (y3628) );
  NAND2x1_ASAP7_75t_R  g7199( .A (n43), .B (n72), .Y (n7207) );
  NAND2x1_ASAP7_75t_R  g7200( .A (n1472), .B (n7207), .Y (y3629) );
  AND3x1_ASAP7_75t_R   g7201( .A (n4129), .B (n3374), .C (n3567), .Y (n7209) );
  NAND2x1_ASAP7_75t_R  g7202( .A (x5), .B (n7209), .Y (y3630) );
  NAND2x1_ASAP7_75t_R  g7203( .A (n12), .B (n3014), .Y (n7211) );
  AND3x1_ASAP7_75t_R   g7204( .A (n7211), .B (n4619), .C (n4618), .Y (y3631) );
  AO21x1_ASAP7_75t_R   g7205( .A1 (n63), .A2 (n363), .B (n530), .Y (y3632) );
  NOR2x1_ASAP7_75t_R   g7206( .A (n12), .B (n403), .Y (n7214) );
  OR3x1_ASAP7_75t_R    g7207( .A (n7214), .B (n529), .C (n29), .Y (y3738) );
  AO21x1_ASAP7_75t_R   g7208( .A1 (n28), .A2 (n388), .B (x3), .Y (n7216) );
  AND2x2_ASAP7_75t_R   g7209( .A (y3738), .B (n7216), .Y (y3634) );
  AND2x2_ASAP7_75t_R   g7210( .A (n6645), .B (n17), .Y (n7218) );
  AO21x1_ASAP7_75t_R   g7211( .A1 (y1467), .A2 (x3), .B (n7218), .Y (y3635) );
  AO21x1_ASAP7_75t_R   g7212( .A1 (n2776), .A2 (n391), .B (n4448), .Y (y3636) );
  AO21x1_ASAP7_75t_R   g7213( .A1 (n2508), .A2 (x1), .B (n1649), .Y (y3637) );
  NOR2x1_ASAP7_75t_R   g7214( .A (n1029), .B (n3433), .Y (y3638) );
  AOI21x1_ASAP7_75t_R  g7215( .A1 (n17), .A2 (n600), .B (n3118), .Y (y3639) );
  AO21x1_ASAP7_75t_R   g7216( .A1 (n17), .A2 (n15), .B (n418), .Y (n7224) );
  AND3x1_ASAP7_75t_R   g7217( .A (n403), .B (x5), .C (x2), .Y (n7225) );
  OR3x1_ASAP7_75t_R    g7218( .A (y2335), .B (n7224), .C (n7225), .Y (n7226) );
  INVx1_ASAP7_75t_R    g7219( .A (n7226), .Y (y3640) );
  OA21x2_ASAP7_75t_R   g7220( .A1 (n139), .A2 (n3376), .B (y3427), .Y (y3641) );
  AO21x1_ASAP7_75t_R   g7221( .A1 (n276), .A2 (x1), .B (y2079), .Y (n7229) );
  AO21x1_ASAP7_75t_R   g7222( .A1 (n129), .A2 (n7229), .B (n2640), .Y (y3642) );
  AO21x1_ASAP7_75t_R   g7223( .A1 (n6610), .A2 (x5), .B (n4541), .Y (y3643) );
  AO21x1_ASAP7_75t_R   g7224( .A1 (n12), .A2 (y2079), .B (y863), .Y (n7232) );
  AOI21x1_ASAP7_75t_R  g7225( .A1 (n7232), .A2 (n2365), .B (n1653), .Y (y3644) );
  OA21x2_ASAP7_75t_R   g7226( .A1 (y3676), .A2 (y1743), .B (n3987), .Y (y3645) );
  INVx1_ASAP7_75t_R    g7227( .A (n3929), .Y (n7235) );
  AND3x1_ASAP7_75t_R   g7228( .A (n7235), .B (y2079), .C (x0), .Y (n7236) );
  INVx1_ASAP7_75t_R    g7229( .A (n7236), .Y (n7237) );
  AO21x1_ASAP7_75t_R   g7230( .A1 (n2718), .A2 (n28), .B (n5250), .Y (y3682) );
  AND2x2_ASAP7_75t_R   g7231( .A (n7237), .B (y3682), .Y (y3646) );
  INVx1_ASAP7_75t_R    g7232( .A (n6792), .Y (n7240) );
  AND3x1_ASAP7_75t_R   g7233( .A (n139), .B (n16), .C (n15), .Y (n7241) );
  OR3x1_ASAP7_75t_R    g7234( .A (n7240), .B (n57), .C (n7241), .Y (y3647) );
  AO21x1_ASAP7_75t_R   g7235( .A1 (n360), .A2 (n3327), .B (n3055), .Y (y3648) );
  AND2x2_ASAP7_75t_R   g7236( .A (n7237), .B (y3427), .Y (y3649) );
  AO21x1_ASAP7_75t_R   g7237( .A1 (n16), .A2 (n2556), .B (n813), .Y (y3650) );
  OA21x2_ASAP7_75t_R   g7238( .A1 (n1137), .A2 (n1431), .B (n4065), .Y (y3651) );
  AO21x1_ASAP7_75t_R   g7239( .A1 (x0), .A2 (x3), .B (x5), .Y (n7247) );
  OA21x2_ASAP7_75t_R   g7240( .A1 (n7247), .A2 (n1110), .B (y3427), .Y (y3652) );
  AO21x1_ASAP7_75t_R   g7241( .A1 (n3646), .A2 (n22), .B (n2994), .Y (n7249) );
  AO32x1_ASAP7_75t_R   g7242( .A1 (n6609), .A2 (n5355), .A3 (y2079), .B1 (x5), .B2 (n7249), .Y (y3653) );
  AND2x2_ASAP7_75t_R   g7243( .A (y1903), .B (n6343), .Y (y3654) );
  AND3x1_ASAP7_75t_R   g7244( .A (n4241), .B (n3143), .C (n632), .Y (y3655) );
  OR3x1_ASAP7_75t_R    g7245( .A (n3112), .B (n6928), .C (n1158), .Y (y3656) );
  OR3x1_ASAP7_75t_R    g7246( .A (n2995), .B (n6928), .C (n1158), .Y (y3657) );
  AO21x1_ASAP7_75t_R   g7247( .A1 (n1246), .A2 (n1247), .B (n462), .Y (y3658) );
  AO21x1_ASAP7_75t_R   g7248( .A1 (y3758), .A2 (x3), .B (n5606), .Y (y3659) );
  AND2x2_ASAP7_75t_R   g7249( .A (n4864), .B (n16), .Y (n7257) );
  NOR2x1_ASAP7_75t_R   g7250( .A (n1208), .B (n7257), .Y (y3660) );
  NOR2x1_ASAP7_75t_R   g7251( .A (n407), .B (n4604), .Y (y3661) );
  NAND2x1_ASAP7_75t_R  g7252( .A (n1163), .B (n388), .Y (n7260) );
  AO21x1_ASAP7_75t_R   g7253( .A1 (n7260), .A2 (x3), .B (n5606), .Y (y3662) );
  AND2x2_ASAP7_75t_R   g7254( .A (n3739), .B (n556), .Y (y3663) );
  AO21x1_ASAP7_75t_R   g7255( .A1 (n22), .A2 (x5), .B (n403), .Y (n7263) );
  OA21x2_ASAP7_75t_R   g7256( .A1 (x0), .A2 (n7263), .B (y1693), .Y (y3664) );
  AND3x1_ASAP7_75t_R   g7257( .A (n290), .B (n360), .C (y2079), .Y (n7265) );
  AO21x1_ASAP7_75t_R   g7258( .A1 (n7235), .A2 (n23), .B (n7265), .Y (y3665) );
  OR3x1_ASAP7_75t_R    g7259( .A (n163), .B (n164), .C (n43), .Y (n7267) );
  NAND2x1_ASAP7_75t_R  g7260( .A (n144), .B (n7267), .Y (y3666) );
  OA21x2_ASAP7_75t_R   g7261( .A1 (n308), .A2 (x3), .B (n3119), .Y (y3667) );
  OA21x2_ASAP7_75t_R   g7262( .A1 (n3519), .A2 (n4117), .B (y2085), .Y (y3668) );
  AND2x2_ASAP7_75t_R   g7263( .A (y1903), .B (n7202), .Y (y3669) );
  NOR2x1_ASAP7_75t_R   g7264( .A (n518), .B (n4719), .Y (y3670) );
  OR3x1_ASAP7_75t_R    g7265( .A (n368), .B (n22), .C (n12), .Y (n7273) );
  INVx1_ASAP7_75t_R    g7266( .A (n7273), .Y (n7274) );
  OR3x1_ASAP7_75t_R    g7267( .A (n7274), .B (n3009), .C (n363), .Y (y3671) );
  AND3x1_ASAP7_75t_R   g7268( .A (n5355), .B (n4907), .C (n388), .Y (n7276) );
  INVx1_ASAP7_75t_R    g7269( .A (n7276), .Y (y3672) );
  AO21x1_ASAP7_75t_R   g7270( .A1 (n495), .A2 (n572), .B (n1190), .Y (n7278) );
  XOR2x2_ASAP7_75t_R   g7271( .A (n7278), .B (x0), .Y (y3673) );
  AND2x2_ASAP7_75t_R   g7272( .A (n572), .B (n3327), .Y (y3674) );
  AND2x2_ASAP7_75t_R   g7273( .A (n3391), .B (y3427), .Y (y3675) );
  OR3x1_ASAP7_75t_R    g7274( .A (n363), .B (n17), .C (x4), .Y (n7282) );
  INVx1_ASAP7_75t_R    g7275( .A (n7282), .Y (n7283) );
  AO21x1_ASAP7_75t_R   g7276( .A1 (n3327), .A2 (x4), .B (n7283), .Y (y3677) );
  OR3x1_ASAP7_75t_R    g7277( .A (n29), .B (n291), .C (n354), .Y (y3678) );
  AO21x1_ASAP7_75t_R   g7278( .A1 (n3138), .A2 (n6220), .B (n45), .Y (y3679) );
  AO32x1_ASAP7_75t_R   g7279( .A1 (n360), .A2 (n3327), .A3 (n310), .B1 (n1158), .B2 (n583), .Y (y3680) );
  AO21x1_ASAP7_75t_R   g7280( .A1 (x0), .A2 (n3474), .B (n4195), .Y (y3681) );
  AND2x2_ASAP7_75t_R   g7281( .A (n1440), .B (n219), .Y (y3683) );
  NAND2x1_ASAP7_75t_R  g7282( .A (n17), .B (n1047), .Y (n7290) );
  AO32x1_ASAP7_75t_R   g7283( .A1 (n17), .A2 (n1047), .A3 (n396), .B1 (y3758), .B2 (n7290), .Y (y3684) );
  AND2x2_ASAP7_75t_R   g7284( .A (n2585), .B (n219), .Y (n7292) );
  AO21x1_ASAP7_75t_R   g7285( .A1 (n17), .A2 (x0), .B (x2), .Y (n7293) );
  OA21x2_ASAP7_75t_R   g7286( .A1 (n7292), .A2 (n15), .B (n7293), .Y (y3685) );
  NAND2x1_ASAP7_75t_R  g7287( .A (x4), .B (n3519), .Y (n7295) );
  AND2x2_ASAP7_75t_R   g7288( .A (n7295), .B (n6866), .Y (y3686) );
  OR3x1_ASAP7_75t_R    g7289( .A (n5410), .B (n1032), .C (x5), .Y (n7297) );
  OA21x2_ASAP7_75t_R   g7290( .A1 (n2994), .A2 (n3426), .B (n7297), .Y (y3687) );
  NAND2x1_ASAP7_75t_R  g7291( .A (x0), .B (n4099), .Y (n7299) );
  AO32x1_ASAP7_75t_R   g7292( .A1 (x0), .A2 (n4099), .A3 (n396), .B1 (y3758), .B2 (n7299), .Y (y3688) );
  AND2x2_ASAP7_75t_R   g7293( .A (y1903), .B (n3648), .Y (y3689) );
  OA21x2_ASAP7_75t_R   g7294( .A1 (n672), .A2 (n5410), .B (y2135), .Y (y3690) );
  AO22x1_ASAP7_75t_R   g7295( .A1 (n22), .A2 (n3004), .B1 (x4), .B2 (n3327), .Y (y3691) );
  AO21x1_ASAP7_75t_R   g7296( .A1 (n997), .A2 (n22), .B (n538), .Y (y3692) );
  AO21x1_ASAP7_75t_R   g7297( .A1 (n3776), .A2 (n3327), .B (n3055), .Y (y3693) );
  AO21x1_ASAP7_75t_R   g7298( .A1 (n1748), .A2 (y2079), .B (n464), .Y (n7306) );
  INVx1_ASAP7_75t_R    g7299( .A (n1114), .Y (n7307) );
  AOI21x1_ASAP7_75t_R  g7300( .A1 (n12), .A2 (n7306), .B (n7307), .Y (y3694) );
  AND3x1_ASAP7_75t_R   g7301( .A (n451), .B (n463), .C (n219), .Y (y3695) );
  AO221x2_ASAP7_75t_R  g7302( .A1 (n1164), .A2 (n4014), .B1 (n4116), .B2 (n1163), .C (n529), .Y (y3696) );
  AND3x1_ASAP7_75t_R   g7303( .A (n1218), .B (n219), .C (n556), .Y (y3697) );
  AND2x2_ASAP7_75t_R   g7304( .A (y1903), .B (n5293), .Y (y3698) );
  AND3x1_ASAP7_75t_R   g7305( .A (n4618), .B (n419), .C (n189), .Y (y3699) );
  OR3x1_ASAP7_75t_R    g7306( .A (n856), .B (n368), .C (x4), .Y (n7314) );
  NAND2x1_ASAP7_75t_R  g7307( .A (n7314), .B (n6551), .Y (y3700) );
  AND2x2_ASAP7_75t_R   g7308( .A (n4755), .B (n189), .Y (y3701) );
  AND2x2_ASAP7_75t_R   g7309( .A (n6871), .B (n189), .Y (y3702) );
  AND2x2_ASAP7_75t_R   g7310( .A (n864), .B (n810), .Y (y3703) );
  AND2x2_ASAP7_75t_R   g7311( .A (n5843), .B (n6343), .Y (y3704) );
  AO21x1_ASAP7_75t_R   g7312( .A1 (n3014), .A2 (n3148), .B (n392), .Y (n7320) );
  NAND2x1_ASAP7_75t_R  g7313( .A (n125), .B (n7320), .Y (y3705) );
  NAND2x1_ASAP7_75t_R  g7314( .A (n16), .B (n2555), .Y (n7322) );
  AO21x1_ASAP7_75t_R   g7315( .A1 (n1424), .A2 (n7322), .B (n195), .Y (y3706) );
  AO21x1_ASAP7_75t_R   g7316( .A1 (n622), .A2 (n418), .B (n3598), .Y (n7324) );
  NOR2x1_ASAP7_75t_R   g7317( .A (n139), .B (n7324), .Y (y3707) );
  NAND2x1_ASAP7_75t_R  g7318( .A (n22), .B (n426), .Y (n7326) );
  AND2x2_ASAP7_75t_R   g7319( .A (n7326), .B (n3261), .Y (y3708) );
  AO21x1_ASAP7_75t_R   g7320( .A1 (n3474), .A2 (x2), .B (n1158), .Y (n7328) );
  XNOR2x2_ASAP7_75t_R  g7321( .A (n5084), .B (n7328), .Y (y3709) );
  AND2x2_ASAP7_75t_R   g7322( .A (n7211), .B (n4618), .Y (y3710) );
  AND2x2_ASAP7_75t_R   g7323( .A (n56), .B (n60), .Y (n7331) );
  AO21x1_ASAP7_75t_R   g7324( .A1 (n7331), .A2 (n17), .B (n4096), .Y (y3711) );
  AND2x2_ASAP7_75t_R   g7325( .A (n917), .B (n1125), .Y (y3712) );
  AO21x1_ASAP7_75t_R   g7326( .A1 (n2718), .A2 (n455), .B (n293), .Y (y3713) );
  AND2x2_ASAP7_75t_R   g7327( .A (n6610), .B (y2079), .Y (y3714) );
  AO21x1_ASAP7_75t_R   g7328( .A1 (n556), .A2 (n3457), .B (n2718), .Y (n7336) );
  AND2x2_ASAP7_75t_R   g7329( .A (n7336), .B (n3797), .Y (y3715) );
  AND3x1_ASAP7_75t_R   g7330( .A (n671), .B (n22), .C (n15), .Y (n7338) );
  INVx1_ASAP7_75t_R    g7331( .A (n7338), .Y (n7339) );
  AND2x2_ASAP7_75t_R   g7332( .A (y2887), .B (n7339), .Y (y3716) );
  OR3x1_ASAP7_75t_R    g7333( .A (n529), .B (n2718), .C (n3009), .Y (y3717) );
  AND2x2_ASAP7_75t_R   g7334( .A (y2085), .B (n6176), .Y (y3718) );
  NOR2x1_ASAP7_75t_R   g7335( .A (n58), .B (n2189), .Y (n7343) );
  NOR2x1_ASAP7_75t_R   g7336( .A (n1245), .B (n7343), .Y (y3719) );
  AO32x1_ASAP7_75t_R   g7337( .A1 (x0), .A2 (n1838), .A3 (n16), .B1 (x1), .B2 (n2557), .Y (y3720) );
  AND2x2_ASAP7_75t_R   g7338( .A (n388), .B (n125), .Y (n7346) );
  NAND2x1_ASAP7_75t_R  g7339( .A (n7346), .B (n5355), .Y (y3721) );
  AO21x1_ASAP7_75t_R   g7340( .A1 (n1572), .A2 (n4459), .B (n3899), .Y (y3722) );
  OR3x1_ASAP7_75t_R    g7341( .A (n7283), .B (n3192), .C (n529), .Y (y3723) );
  AND2x2_ASAP7_75t_R   g7342( .A (n3794), .B (n3316), .Y (n7350) );
  AO21x1_ASAP7_75t_R   g7343( .A1 (n1572), .A2 (n4459), .B (n7350), .Y (y3724) );
  AND3x1_ASAP7_75t_R   g7344( .A (y3852), .B (n352), .C (n17), .Y (n7352) );
  OR3x1_ASAP7_75t_R    g7345( .A (n7283), .B (n7352), .C (n529), .Y (y3725) );
  AO21x1_ASAP7_75t_R   g7346( .A1 (n3148), .A2 (n2776), .B (n7197), .Y (y3726) );
  AO21x1_ASAP7_75t_R   g7347( .A1 (x0), .A2 (x1), .B (n22), .Y (n7355) );
  AO21x1_ASAP7_75t_R   g7348( .A1 (y2079), .A2 (n7355), .B (n1150), .Y (y3727) );
  OR3x1_ASAP7_75t_R    g7349( .A (n529), .B (n1158), .C (n3192), .Y (y3728) );
  OR3x1_ASAP7_75t_R    g7350( .A (n7352), .B (n1158), .C (n529), .Y (y3729) );
  AO21x1_ASAP7_75t_R   g7351( .A1 (n12), .A2 (n4739), .B (y2916), .Y (y3730) );
  AND2x2_ASAP7_75t_R   g7352( .A (y1903), .B (n455), .Y (y3731) );
  AO21x1_ASAP7_75t_R   g7353( .A1 (x5), .A2 (x3), .B (n22), .Y (n7361) );
  AO21x1_ASAP7_75t_R   g7354( .A1 (y2079), .A2 (n17), .B (x4), .Y (n7362) );
  NAND2x1_ASAP7_75t_R  g7355( .A (n7361), .B (n7362), .Y (y3799) );
  AND2x2_ASAP7_75t_R   g7356( .A (y3799), .B (x0), .Y (y3733) );
  AND2x2_ASAP7_75t_R   g7357( .A (y1903), .B (n451), .Y (y3734) );
  AND2x2_ASAP7_75t_R   g7358( .A (y1903), .B (n2797), .Y (y3735) );
  AO21x1_ASAP7_75t_R   g7359( .A1 (n3736), .A2 (n3327), .B (n29), .Y (y3736) );
  AO21x1_ASAP7_75t_R   g7360( .A1 (n5819), .A2 (y2079), .B (n6821), .Y (y3737) );
  AND2x2_ASAP7_75t_R   g7361( .A (n980), .B (n387), .Y (y3739) );
  AND2x2_ASAP7_75t_R   g7362( .A (y1903), .B (n632), .Y (y3740) );
  OR3x1_ASAP7_75t_R    g7363( .A (y3758), .B (n2718), .C (n1158), .Y (y3741) );
  OA21x2_ASAP7_75t_R   g7364( .A1 (x1), .A2 (n3417), .B (n1272), .Y (y3742) );
  AND2x2_ASAP7_75t_R   g7365( .A (n4824), .B (n419), .Y (y3743) );
  AO21x1_ASAP7_75t_R   g7366( .A1 (n15), .A2 (n22), .B (x3), .Y (n7374) );
  AND2x2_ASAP7_75t_R   g7367( .A (n360), .B (n7374), .Y (n7375) );
  AO21x1_ASAP7_75t_R   g7368( .A1 (n7375), .A2 (y2079), .B (n2050), .Y (y3744) );
  OA22x2_ASAP7_75t_R   g7369( .A1 (n291), .A2 (n5419), .B1 (y2068), .B2 (n15), .Y (y3745) );
  AO21x1_ASAP7_75t_R   g7370( .A1 (n360), .A2 (n3267), .B (x5), .Y (n7378) );
  AND2x2_ASAP7_75t_R   g7371( .A (n6460), .B (n7378), .Y (y3746) );
  OR3x1_ASAP7_75t_R    g7372( .A (n2999), .B (n403), .C (x5), .Y (n7380) );
  OA21x2_ASAP7_75t_R   g7373( .A1 (n378), .A2 (y2079), .B (n7380), .Y (y3747) );
  NOR2x1_ASAP7_75t_R   g7374( .A (n2897), .B (n1462), .Y (y3748) );
  INVx1_ASAP7_75t_R    g7375( .A (n1782), .Y (n7383) );
  NOR2x1_ASAP7_75t_R   g7376( .A (n1339), .B (n7383), .Y (y3749) );
  AND2x2_ASAP7_75t_R   g7377( .A (n1110), .B (n3005), .Y (y3750) );
  AO21x1_ASAP7_75t_R   g7378( .A1 (n556), .A2 (x3), .B (n6928), .Y (y3751) );
  AND2x2_ASAP7_75t_R   g7379( .A (n1620), .B (n5575), .Y (y3752) );
  OR3x1_ASAP7_75t_R    g7380( .A (n296), .B (n297), .C (n5679), .Y (y3753) );
  AO21x1_ASAP7_75t_R   g7381( .A1 (n291), .A2 (n740), .B (n293), .Y (y3755) );
  AO21x1_ASAP7_75t_R   g7382( .A1 (n546), .A2 (n463), .B (x0), .Y (y3756) );
  AND2x2_ASAP7_75t_R   g7383( .A (n5932), .B (n3119), .Y (y3757) );
  NOR2x1_ASAP7_75t_R   g7384( .A (x5), .B (n4535), .Y (n7392) );
  AO21x1_ASAP7_75t_R   g7385( .A1 (n7235), .A2 (x5), .B (n7392), .Y (y3759) );
  AND2x2_ASAP7_75t_R   g7386( .A (y3132), .B (n6566), .Y (y3760) );
  NOR2x1_ASAP7_75t_R   g7387( .A (n352), .B (n63), .Y (n7395) );
  NOR2x1_ASAP7_75t_R   g7388( .A (n4192), .B (n7395), .Y (y3761) );
  AO21x1_ASAP7_75t_R   g7389( .A1 (y863), .A2 (x2), .B (n17), .Y (n7397) );
  OA21x2_ASAP7_75t_R   g7390( .A1 (n2873), .A2 (x3), .B (n7397), .Y (y3762) );
  AND2x2_ASAP7_75t_R   g7391( .A (n3325), .B (y2079), .Y (n7399) );
  AO21x1_ASAP7_75t_R   g7392( .A1 (n22), .A2 (n397), .B (n7399), .Y (y3763) );
  AND2x2_ASAP7_75t_R   g7393( .A (n6566), .B (n367), .Y (y3764) );
  AND2x2_ASAP7_75t_R   g7394( .A (y3615), .B (n419), .Y (y3765) );
  INVx1_ASAP7_75t_R    g7395( .A (n5081), .Y (n7403) );
  AO21x1_ASAP7_75t_R   g7396( .A1 (n3457), .A2 (n2246), .B (n7403), .Y (y3766) );
  AO21x1_ASAP7_75t_R   g7397( .A1 (n1305), .A2 (n1743), .B (n1745), .Y (y3767) );
  AO21x1_ASAP7_75t_R   g7398( .A1 (n660), .A2 (n406), .B (x0), .Y (n7406) );
  OA21x2_ASAP7_75t_R   g7399( .A1 (y1260), .A2 (n12), .B (n7406), .Y (y3768) );
  NOR2x1_ASAP7_75t_R   g7400( .A (n3118), .B (n921), .Y (y3769) );
  NOR2x1_ASAP7_75t_R   g7401( .A (x5), .B (n3883), .Y (n7409) );
  AO21x1_ASAP7_75t_R   g7402( .A1 (n7235), .A2 (x5), .B (n7409), .Y (y3770) );
  AO21x1_ASAP7_75t_R   g7403( .A1 (n137), .A2 (x5), .B (n4844), .Y (n7411) );
  AO21x1_ASAP7_75t_R   g7404( .A1 (n137), .A2 (y2079), .B (n3284), .Y (n7412) );
  AND2x2_ASAP7_75t_R   g7405( .A (n7411), .B (n7412), .Y (y3771) );
  NOR2x1_ASAP7_75t_R   g7406( .A (n518), .B (n231), .Y (n7414) );
  AND3x1_ASAP7_75t_R   g7407( .A (n58), .B (n22), .C (n16), .Y (n7415) );
  INVx1_ASAP7_75t_R    g7408( .A (n7415), .Y (n7416) );
  OA21x2_ASAP7_75t_R   g7409( .A1 (x0), .A2 (n7414), .B (n7416), .Y (y3772) );
  INVx1_ASAP7_75t_R    g7410( .A (n4844), .Y (n7418) );
  AO32x1_ASAP7_75t_R   g7411( .A1 (n2966), .A2 (x4), .A3 (n1062), .B1 (n672), .B2 (n7418), .Y (y3773) );
  OA21x2_ASAP7_75t_R   g7412( .A1 (n434), .A2 (n1942), .B (n935), .Y (y3774) );
  AO21x1_ASAP7_75t_R   g7413( .A1 (n3567), .A2 (x3), .B (n3659), .Y (n7421) );
  OR3x1_ASAP7_75t_R    g7414( .A (n7421), .B (n3637), .C (x5), .Y (n7422) );
  INVx1_ASAP7_75t_R    g7415( .A (n5127), .Y (n7423) );
  OR3x1_ASAP7_75t_R    g7416( .A (n291), .B (n7423), .C (y2079), .Y (y3790) );
  AND2x2_ASAP7_75t_R   g7417( .A (n7422), .B (y3790), .Y (y3775) );
  OR3x1_ASAP7_75t_R    g7418( .A (n1004), .B (n1778), .C (n527), .Y (y3776) );
  AO21x1_ASAP7_75t_R   g7419( .A1 (n360), .A2 (n290), .B (n740), .Y (n7427) );
  AO21x1_ASAP7_75t_R   g7420( .A1 (n137), .A2 (n22), .B (n3474), .Y (n7428) );
  AND2x2_ASAP7_75t_R   g7421( .A (n7427), .B (n7428), .Y (y3777) );
  AND3x1_ASAP7_75t_R   g7422( .A (n556), .B (n3457), .C (x2), .Y (n7430) );
  AO21x1_ASAP7_75t_R   g7423( .A1 (n4755), .A2 (n3297), .B (n7430), .Y (y3778) );
  AND3x1_ASAP7_75t_R   g7424( .A (n1300), .B (n137), .C (n72), .Y (n7432) );
  AO21x1_ASAP7_75t_R   g7425( .A1 (n218), .A2 (n1299), .B (n7432), .Y (n7433) );
  OR3x1_ASAP7_75t_R    g7426( .A (n7433), .B (n130), .C (n13), .Y (y3779) );
  AO21x1_ASAP7_75t_R   g7427( .A1 (n3567), .A2 (x5), .B (n3374), .Y (n7435) );
  AND2x2_ASAP7_75t_R   g7428( .A (n7435), .B (n3119), .Y (y3780) );
  OA21x2_ASAP7_75t_R   g7429( .A1 (n856), .A2 (n3777), .B (n5178), .Y (y3781) );
  NAND2x1_ASAP7_75t_R  g7430( .A (n5127), .B (n290), .Y (n7438) );
  AO21x1_ASAP7_75t_R   g7431( .A1 (n7438), .A2 (n1265), .B (n349), .Y (y3782) );
  OA21x2_ASAP7_75t_R   g7432( .A1 (n1339), .A2 (n1424), .B (n2915), .Y (y3783) );
  OR3x1_ASAP7_75t_R    g7433( .A (y3758), .B (n163), .C (n164), .Y (y3784) );
  INVx1_ASAP7_75t_R    g7434( .A (n3227), .Y (n7442) );
  OA21x2_ASAP7_75t_R   g7435( .A1 (n164), .A2 (n406), .B (n7442), .Y (y3785) );
  AND2x2_ASAP7_75t_R   g7436( .A (y1693), .B (n3143), .Y (n7444) );
  AO21x1_ASAP7_75t_R   g7437( .A1 (n639), .A2 (n3144), .B (n7444), .Y (y3786) );
  AO21x1_ASAP7_75t_R   g7438( .A1 (y2632), .A2 (n4935), .B (y863), .Y (y3787) );
  AO21x1_ASAP7_75t_R   g7439( .A1 (y2079), .A2 (x2), .B (n518), .Y (n7447) );
  INVx1_ASAP7_75t_R    g7440( .A (n7447), .Y (n7448) );
  AO21x1_ASAP7_75t_R   g7441( .A1 (n7448), .A2 (n3000), .B (x3), .Y (n7449) );
  NAND2x1_ASAP7_75t_R  g7442( .A (n292), .B (n7449), .Y (y3788) );
  AO21x1_ASAP7_75t_R   g7443( .A1 (n16), .A2 (n22), .B (n363), .Y (n7451) );
  AO21x1_ASAP7_75t_R   g7444( .A1 (n143), .A2 (n455), .B (n7451), .Y (y3789) );
  NAND2x1_ASAP7_75t_R  g7445( .A (n976), .B (n312), .Y (y3791) );
  INVx1_ASAP7_75t_R    g7446( .A (n7247), .Y (n7454) );
  NAND2x1_ASAP7_75t_R  g7447( .A (n3370), .B (n7454), .Y (n7455) );
  AND2x2_ASAP7_75t_R   g7448( .A (n7455), .B (n3475), .Y (y3792) );
  NAND2x1_ASAP7_75t_R  g7449( .A (y2079), .B (n328), .Y (n7457) );
  AO21x1_ASAP7_75t_R   g7450( .A1 (n382), .A2 (n681), .B (y2079), .Y (y3797) );
  OA21x2_ASAP7_75t_R   g7451( .A1 (n7457), .A2 (n3039), .B (y3797), .Y (y3793) );
  AO21x1_ASAP7_75t_R   g7452( .A1 (y2079), .A2 (n3482), .B (n638), .Y (y3794) );
  INVx1_ASAP7_75t_R    g7453( .A (n391), .Y (n7461) );
  AO32x1_ASAP7_75t_R   g7454( .A1 (y3293), .A2 (n125), .A3 (n391), .B1 (n7461), .B2 (n429), .Y (y3795) );
  OR3x1_ASAP7_75t_R    g7455( .A (n4908), .B (n3009), .C (n529), .Y (y3796) );
  OA21x2_ASAP7_75t_R   g7456( .A1 (n2226), .A2 (n143), .B (n1640), .Y (y3798) );
  AO21x1_ASAP7_75t_R   g7457( .A1 (n3327), .A2 (x4), .B (n3055), .Y (y3800) );
  OR3x1_ASAP7_75t_R    g7458( .A (n1158), .B (n421), .C (n5385), .Y (y3801) );
  NAND2x1_ASAP7_75t_R  g7459( .A (n4708), .B (n360), .Y (n7467) );
  INVx1_ASAP7_75t_R    g7460( .A (n7467), .Y (n7468) );
  AO32x1_ASAP7_75t_R   g7461( .A1 (n15), .A2 (n455), .A3 (n7468), .B1 (n7467), .B2 (n5090), .Y (y3803) );
  INVx1_ASAP7_75t_R    g7462( .A (n356), .Y (n7470) );
  OR3x1_ASAP7_75t_R    g7463( .A (n291), .B (n29), .C (n7470), .Y (y3804) );
  NOR2x1_ASAP7_75t_R   g7464( .A (n111), .B (n1613), .Y (y3805) );
  AND2x2_ASAP7_75t_R   g7465( .A (n1891), .B (y1958), .Y (y3806) );
  AND2x2_ASAP7_75t_R   g7466( .A (n415), .B (y2079), .Y (n7474) );
  OR3x1_ASAP7_75t_R    g7467( .A (n3055), .B (n2994), .C (n7474), .Y (y3807) );
  AO21x1_ASAP7_75t_R   g7468( .A1 (n466), .A2 (n1093), .B (n972), .Y (y3809) );
  AO21x1_ASAP7_75t_R   g7469( .A1 (n604), .A2 (n994), .B (n3450), .Y (y3810) );
  AND2x2_ASAP7_75t_R   g7470( .A (n3966), .B (n1383), .Y (y3811) );
  AO21x1_ASAP7_75t_R   g7471( .A1 (n455), .A2 (n84), .B (n2718), .Y (n7479) );
  AO21x1_ASAP7_75t_R   g7472( .A1 (n7479), .A2 (n556), .B (n4403), .Y (y3812) );
  OR3x1_ASAP7_75t_R    g7473( .A (n392), .B (n15), .C (x3), .Y (n7481) );
  AND2x2_ASAP7_75t_R   g7474( .A (n7481), .B (n4618), .Y (y3813) );
  AND3x1_ASAP7_75t_R   g7475( .A (n1062), .B (n388), .C (n28), .Y (n7483) );
  AO21x1_ASAP7_75t_R   g7476( .A1 (n1838), .A2 (n419), .B (n7483), .Y (n7484) );
  NOR2x1_ASAP7_75t_R   g7477( .A (y2079), .B (n4647), .Y (n7485) );
  INVx1_ASAP7_75t_R    g7478( .A (n7485), .Y (n7486) );
  NAND2x1_ASAP7_75t_R  g7479( .A (n7484), .B (n7486), .Y (y3814) );
  AO21x1_ASAP7_75t_R   g7480( .A1 (x3), .A2 (n3027), .B (n337), .Y (n7488) );
  AO21x1_ASAP7_75t_R   g7481( .A1 (x5), .A2 (n3143), .B (n7488), .Y (n7489) );
  AO21x1_ASAP7_75t_R   g7482( .A1 (n4374), .A2 (n401), .B (y2079), .Y (n7490) );
  AND2x2_ASAP7_75t_R   g7483( .A (n7489), .B (n7490), .Y (y3815) );
  AO21x1_ASAP7_75t_R   g7484( .A1 (y2079), .A2 (n1175), .B (n1150), .Y (y3816) );
  AO21x1_ASAP7_75t_R   g7485( .A1 (y3758), .A2 (x2), .B (n6572), .Y (y3817) );
  INVx1_ASAP7_75t_R    g7486( .A (n3361), .Y (n7494) );
  OA211x2_ASAP7_75t_R  g7487( .A1 (n396), .A2 (n76), .B (n1572), .C (n7494), .Y (y3818) );
  _const1_             g7488( .z (y3819) );
  AND2x2_ASAP7_75t_R   g7489( .A (y3615), .B (n5224), .Y (y3820) );
  OR3x1_ASAP7_75t_R    g7490( .A (n184), .B (n271), .C (n262), .Y (y3821) );
  AO21x1_ASAP7_75t_R   g7491( .A1 (n1047), .A2 (x1), .B (n1095), .Y (y3822) );
  AO21x1_ASAP7_75t_R   g7492( .A1 (n17), .A2 (n6291), .B (n164), .Y (n7500) );
  INVx1_ASAP7_75t_R    g7493( .A (n7500), .Y (n7501) );
  AO32x1_ASAP7_75t_R   g7494( .A1 (n388), .A2 (n28), .A3 (n7500), .B1 (n7501), .B2 (y3758), .Y (y3823) );
  NAND2x1_ASAP7_75t_R  g7495( .A (x5), .B (n5174), .Y (y3844) );
  OA21x2_ASAP7_75t_R   g7496( .A1 (x5), .A2 (n5174), .B (y3844), .Y (y3824) );
  INVx1_ASAP7_75t_R    g7497( .A (n3617), .Y (n7505) );
  AO21x1_ASAP7_75t_R   g7498( .A1 (n556), .A2 (x2), .B (n3617), .Y (n7506) );
  AO32x1_ASAP7_75t_R   g7499( .A1 (n7505), .A2 (n291), .A3 (n3297), .B1 (x3), .B2 (n7506), .Y (y3825) );
  XOR2x2_ASAP7_75t_R   g7500( .A (n6387), .B (y2079), .Y (y3826) );
  AO21x1_ASAP7_75t_R   g7501( .A1 (n15), .A2 (n4903), .B (n421), .Y (n7509) );
  XOR2x2_ASAP7_75t_R   g7502( .A (n7509), .B (n6272), .Y (y3827) );
  AO21x1_ASAP7_75t_R   g7503( .A1 (n144), .A2 (n81), .B (n4291), .Y (y3828) );
  AO21x1_ASAP7_75t_R   g7504( .A1 (n6176), .A2 (n366), .B (n218), .Y (y3829) );
  AND2x2_ASAP7_75t_R   g7505( .A (y2610), .B (n6733), .Y (y3830) );
  AO21x1_ASAP7_75t_R   g7506( .A1 (n3804), .A2 (y2079), .B (n76), .Y (n7514) );
  AO21x1_ASAP7_75t_R   g7507( .A1 (n5910), .A2 (n7514), .B (n7485), .Y (y3832) );
  AO21x1_ASAP7_75t_R   g7508( .A1 (n64), .A2 (n63), .B (x3), .Y (n7516) );
  NAND2x1_ASAP7_75t_R  g7509( .A (n7516), .B (n2594), .Y (y3833) );
  NOR2x1_ASAP7_75t_R   g7510( .A (n4150), .B (n4983), .Y (y3834) );
  AO21x1_ASAP7_75t_R   g7511( .A1 (x2), .A2 (n17), .B (n90), .Y (n7519) );
  AND3x1_ASAP7_75t_R   g7512( .A (n4261), .B (n7519), .C (n244), .Y (y3835) );
  AO21x1_ASAP7_75t_R   g7513( .A1 (n319), .A2 (n22), .B (n3285), .Y (n7521) );
  AND2x2_ASAP7_75t_R   g7514( .A (n5297), .B (n7521), .Y (y3836) );
  NAND2x1_ASAP7_75t_R  g7515( .A (n15), .B (n647), .Y (n7523) );
  OR3x1_ASAP7_75t_R    g7516( .A (n291), .B (n15), .C (n293), .Y (n7524) );
  OA21x2_ASAP7_75t_R   g7517( .A1 (n5827), .A2 (n7523), .B (n7524), .Y (y3837) );
  AND3x1_ASAP7_75t_R   g7518( .A (n17), .B (x0), .C (x1), .Y (n7526) );
  INVx1_ASAP7_75t_R    g7519( .A (n7526), .Y (n7527) );
  INVx1_ASAP7_75t_R    g7520( .A (n5393), .Y (n7528) );
  OA21x2_ASAP7_75t_R   g7521( .A1 (n7528), .A2 (n7526), .B (n228), .Y (n7529) );
  AO32x1_ASAP7_75t_R   g7522( .A1 (x2), .A2 (n7527), .A3 (n5393), .B1 (n7529), .B2 (n15), .Y (y3838) );
  AO21x1_ASAP7_75t_R   g7523( .A1 (y9), .A2 (n890), .B (n2880), .Y (y3839) );
  AO21x1_ASAP7_75t_R   g7524( .A1 (n97), .A2 (x3), .B (n3294), .Y (n7532) );
  OA211x2_ASAP7_75t_R  g7525( .A1 (n7532), .A2 (n22), .B (n740), .C (n4109), .Y (n7533) );
  INVx1_ASAP7_75t_R    g7526( .A (n7533), .Y (y3840) );
  INVx1_ASAP7_75t_R    g7527( .A (n3524), .Y (n7535) );
  AO21x1_ASAP7_75t_R   g7528( .A1 (x2), .A2 (x4), .B (y2079), .Y (n7536) );
  INVx1_ASAP7_75t_R    g7529( .A (n7536), .Y (n7537) );
  OA33x2_ASAP7_75t_R   g7530( .A1 (n211), .A2 (y2079), .A3 (n7535), .B1 (n3618), .B2 (n1269), .B3 (n7537), .Y (y3841) );
  AND2x2_ASAP7_75t_R   g7531( .A (n3762), .B (n366), .Y (n7539) );
  AO21x1_ASAP7_75t_R   g7532( .A1 (n3493), .A2 (x4), .B (n7539), .Y (y3842) );
  AND2x2_ASAP7_75t_R   g7533( .A (n3898), .B (n4090), .Y (y3843) );
  OA21x2_ASAP7_75t_R   g7534( .A1 (n2959), .A2 (n1643), .B (n1066), .Y (y3845) );
  NAND2x1_ASAP7_75t_R  g7535( .A (y2079), .B (n4107), .Y (n7543) );
  AO21x1_ASAP7_75t_R   g7536( .A1 (y2079), .A2 (n4107), .B (n29), .Y (n7544) );
  AO32x1_ASAP7_75t_R   g7537( .A1 (n28), .A2 (n7543), .A3 (n217), .B1 (n218), .B2 (n7544), .Y (n7545) );
  INVx1_ASAP7_75t_R    g7538( .A (n7545), .Y (y3846) );
  INVx1_ASAP7_75t_R    g7539( .A (n6220), .Y (n7547) );
  OR3x1_ASAP7_75t_R    g7540( .A (n7547), .B (n4340), .C (x3), .Y (n7548) );
  AO21x1_ASAP7_75t_R   g7541( .A1 (n4341), .A2 (n4528), .B (n17), .Y (n7549) );
  AND2x2_ASAP7_75t_R   g7542( .A (n7548), .B (n7549), .Y (y3847) );
  AO21x1_ASAP7_75t_R   g7543( .A1 (n455), .A2 (n76), .B (n81), .Y (n7551) );
  AOI21x1_ASAP7_75t_R  g7544( .A1 (n7551), .A2 (n396), .B (y2771), .Y (y3848) );
  AO21x1_ASAP7_75t_R   g7545( .A1 (n46), .A2 (n47), .B (n143), .Y (y3849) );
  AO21x1_ASAP7_75t_R   g7546( .A1 (n301), .A2 (n299), .B (x3), .Y (n7554) );
  AND2x2_ASAP7_75t_R   g7547( .A (n7554), .B (n3882), .Y (y3850) );
  NAND2x1_ASAP7_75t_R  g7548( .A (x3), .B (n5256), .Y (n7556) );
  AO32x1_ASAP7_75t_R   g7549( .A1 (x3), .A2 (n5256), .A3 (n4551), .B1 (n4550), .B2 (n7556), .Y (y3851) );
  NOR2x1_ASAP7_75t_R   g7550( .A (n3494), .B (n4983), .Y (y3853) );
  AO32x1_ASAP7_75t_R   g7551( .A1 (n5094), .A2 (n3828), .A3 (x4), .B1 (n3944), .B2 (n7532), .Y (y3854) );
  OA21x2_ASAP7_75t_R   g7552( .A1 (n1190), .A2 (y195), .B (n3879), .Y (y3855) );
  NAND2x1_ASAP7_75t_R  g7553( .A (n137), .B (n6322), .Y (n7561) );
  AO21x1_ASAP7_75t_R   g7554( .A1 (n97), .A2 (x3), .B (n4107), .Y (n7562) );
  OA21x2_ASAP7_75t_R   g7555( .A1 (n7561), .A2 (n3907), .B (n7562), .Y (y3856) );
  OR3x1_ASAP7_75t_R    g7556( .A (n1184), .B (n43), .C (n529), .Y (y3857) );
  AND3x1_ASAP7_75t_R   g7557( .A (n5072), .B (n3469), .C (n3567), .Y (n7565) );
  AO21x1_ASAP7_75t_R   g7558( .A1 (n4551), .A2 (n3638), .B (n7565), .Y (n7566) );
  AO21x1_ASAP7_75t_R   g7559( .A1 (x2), .A2 (y2079), .B (n7566), .Y (y3858) );
  INVx1_ASAP7_75t_R    g7560( .A (n7561), .Y (n7568) );
  AO221x2_ASAP7_75t_R  g7561( .A1 (n7568), .A2 (n22), .B1 (x4), .B2 (n7561), .C (n6390), .Y (y3859) );
  AO21x1_ASAP7_75t_R   g7562( .A1 (n3133), .A2 (n455), .B (n3135), .Y (y3860) );
  NOR2x1_ASAP7_75t_R   g7563( .A (n366), .B (n4972), .Y (n7571) );
  NOR2x1_ASAP7_75t_R   g7564( .A (n7571), .B (n5451), .Y (y3861) );
  OA21x2_ASAP7_75t_R   g7565( .A1 (n217), .A2 (n28), .B (n4090), .Y (y3862) );
  AO32x1_ASAP7_75t_R   g7566( .A1 (n4216), .A2 (x4), .A3 (n72), .B1 (n3316), .B2 (n4727), .Y (n7574) );
  NAND2x1_ASAP7_75t_R  g7567( .A (n3794), .B (n7574), .Y (y3863) );
  AO32x1_ASAP7_75t_R   g7568( .A1 (n144), .A2 (n1954), .A3 (n15), .B1 (x2), .B2 (y1356), .Y (y3864) );
  OR3x1_ASAP7_75t_R    g7569( .A (n4648), .B (y2079), .C (n3992), .Y (y3865) );
  OR3x1_ASAP7_75t_R    g7570( .A (n4483), .B (n3628), .C (n2999), .Y (y3866) );
  AO21x1_ASAP7_75t_R   g7571( .A1 (x5), .A2 (n2989), .B (n4841), .Y (y3867) );
  AND3x1_ASAP7_75t_R   g7572( .A (y1903), .B (n3648), .C (n84), .Y (y3868) );
  AO21x1_ASAP7_75t_R   g7573( .A1 (n17), .A2 (x2), .B (y2466), .Y (n7581) );
  AO21x1_ASAP7_75t_R   g7574( .A1 (x2), .A2 (n556), .B (n7581), .Y (n7582) );
  AO21x1_ASAP7_75t_R   g7575( .A1 (x3), .A2 (n3617), .B (n7582), .Y (y3869) );
  OA21x2_ASAP7_75t_R   g7576( .A1 (x5), .A2 (n3311), .B (y2296), .Y (y3870) );
  AO21x1_ASAP7_75t_R   g7577( .A1 (n382), .A2 (n97), .B (n1269), .Y (n7585) );
  AO21x1_ASAP7_75t_R   g7578( .A1 (x4), .A2 (n5996), .B (n7585), .Y (y3871) );
  OA21x2_ASAP7_75t_R   g7579( .A1 (n3033), .A2 (n3035), .B (n2254), .Y (y3872) );
  INVx1_ASAP7_75t_R    g7580( .A (n3565), .Y (n7588) );
  AND2x2_ASAP7_75t_R   g7581( .A (x5), .B (x2), .Y (n7589) );
  OR3x1_ASAP7_75t_R    g7582( .A (n7589), .B (n22), .C (n17), .Y (n7590) );
  INVx1_ASAP7_75t_R    g7583( .A (n7590), .Y (n7591) );
  AO21x1_ASAP7_75t_R   g7584( .A1 (x2), .A2 (n7588), .B (n7591), .Y (y3873) );
  AO21x1_ASAP7_75t_R   g7585( .A1 (n243), .A2 (n15), .B (x0), .Y (n7593) );
  AND2x2_ASAP7_75t_R   g7586( .A (n2358), .B (n7593), .Y (y3874) );
  OA21x2_ASAP7_75t_R   g7587( .A1 (x5), .A2 (n4581), .B (y2737), .Y (y3875) );
  OR3x1_ASAP7_75t_R    g7588( .A (x5), .B (x3), .C (x2), .Y (n7596) );
  INVx1_ASAP7_75t_R    g7589( .A (n7596), .Y (n7597) );
  OA211x2_ASAP7_75t_R  g7590( .A1 (n7597), .A2 (n7589), .B (n5666), .C (x4), .Y (n7598) );
  INVx1_ASAP7_75t_R    g7591( .A (n5666), .Y (n7599) );
  INVx1_ASAP7_75t_R    g7592( .A (n7589), .Y (n7600) );
  OA211x2_ASAP7_75t_R  g7593( .A1 (n7599), .A2 (n22), .B (n7600), .C (n7596), .Y (n7601) );
  NOR2x1_ASAP7_75t_R   g7594( .A (n7598), .B (n7601), .Y (y3876) );
  NOR2x1_ASAP7_75t_R   g7595( .A (n3338), .B (n3237), .Y (n7603) );
  INVx1_ASAP7_75t_R    g7596( .A (n7603), .Y (n7604) );
  AO21x1_ASAP7_75t_R   g7597( .A1 (n28), .A2 (n290), .B (n756), .Y (n7605) );
  AND2x2_ASAP7_75t_R   g7598( .A (n7604), .B (n7605), .Y (y3877) );
  AO21x1_ASAP7_75t_R   g7599( .A1 (n76), .A2 (n228), .B (n2922), .Y (y3878) );
  AO21x1_ASAP7_75t_R   g7600( .A1 (n2246), .A2 (n3457), .B (n2994), .Y (y3879) );
  AO21x1_ASAP7_75t_R   g7601( .A1 (n660), .A2 (x2), .B (n6043), .Y (n7609) );
  AND2x2_ASAP7_75t_R   g7602( .A (n7609), .B (n3282), .Y (y3880) );
  NOR2x1_ASAP7_75t_R   g7603( .A (n671), .B (n3144), .Y (n7611) );
  AND2x2_ASAP7_75t_R   g7604( .A (n4241), .B (n7611), .Y (y3881) );
  AO32x1_ASAP7_75t_R   g7605( .A1 (n137), .A2 (n5108), .A3 (n72), .B1 (n4089), .B2 (n4102), .Y (y3882) );
  AO21x1_ASAP7_75t_R   g7606( .A1 (y1378), .A2 (x1), .B (n3050), .Y (y3884) );
  OA21x2_ASAP7_75t_R   g7607( .A1 (n421), .A2 (n3000), .B (n3302), .Y (n7615) );
  XOR2x2_ASAP7_75t_R   g7608( .A (n7615), .B (n17), .Y (y3885) );
  OR3x1_ASAP7_75t_R    g7609( .A (n276), .B (x5), .C (x1), .Y (n7617) );
  NAND2x1_ASAP7_75t_R  g7610( .A (n7617), .B (n1291), .Y (y3886) );
  NAND2x1_ASAP7_75t_R  g7611( .A (x5), .B (n5116), .Y (n7619) );
  AO21x1_ASAP7_75t_R   g7612( .A1 (n4643), .A2 (n7619), .B (n3310), .Y (y3887) );
  AND3x1_ASAP7_75t_R   g7613( .A (n97), .B (n740), .C (n17), .Y (n7621) );
  OR3x1_ASAP7_75t_R    g7614( .A (n3719), .B (n7621), .C (n3568), .Y (y3888) );
  AND2x2_ASAP7_75t_R   g7615( .A (n3024), .B (y2079), .Y (n7623) );
  AO21x1_ASAP7_75t_R   g7616( .A1 (n22), .A2 (n3828), .B (n7623), .Y (y3889) );
  AO21x1_ASAP7_75t_R   g7617( .A1 (x5), .A2 (n17), .B (n3028), .Y (n7625) );
  AO21x1_ASAP7_75t_R   g7618( .A1 (n3286), .A2 (n7625), .B (n628), .Y (y3890) );
  AND2x2_ASAP7_75t_R   g7619( .A (n2748), .B (x0), .Y (n7627) );
  AO21x1_ASAP7_75t_R   g7620( .A1 (x0), .A2 (n17), .B (n64), .Y (n7628) );
  OA21x2_ASAP7_75t_R   g7621( .A1 (n7627), .A2 (n2556), .B (n7628), .Y (y3891) );
  AND2x2_ASAP7_75t_R   g7622( .A (n3391), .B (y2085), .Y (y3892) );
  AND3x1_ASAP7_75t_R   g7623( .A (n756), .B (x3), .C (x4), .Y (n7631) );
  NOR2x1_ASAP7_75t_R   g7624( .A (n4279), .B (n7631), .Y (y3893) );
  AND2x2_ASAP7_75t_R   g7625( .A (n5243), .B (y2079), .Y (n7633) );
  OR3x1_ASAP7_75t_R    g7626( .A (n7633), .B (n5117), .C (n3310), .Y (y3894) );
  AO22x1_ASAP7_75t_R   g7627( .A1 (n6190), .A2 (x2), .B1 (n3183), .B2 (x3), .Y (y3895) );
  AO21x1_ASAP7_75t_R   g7628( .A1 (y2079), .A2 (n84), .B (y3800), .Y (y3896) );
  AO21x1_ASAP7_75t_R   g7629( .A1 (x5), .A2 (n5117), .B (n286), .Y (n7637) );
  AO21x1_ASAP7_75t_R   g7630( .A1 (n15), .A2 (n287), .B (n7637), .Y (y3897) );
  AO21x1_ASAP7_75t_R   g7631( .A1 (n2980), .A2 (n4821), .B (n286), .Y (y3898) );
  AO21x1_ASAP7_75t_R   g7632( .A1 (x1), .A2 (n58), .B (n4627), .Y (y3899) );
  AO32x1_ASAP7_75t_R   g7633( .A1 (n312), .A2 (x0), .A3 (n466), .B1 (x4), .B2 (n6401), .Y (y3900) );
  AO21x1_ASAP7_75t_R   g7634( .A1 (y2079), .A2 (n228), .B (n3732), .Y (n7642) );
  AND2x2_ASAP7_75t_R   g7635( .A (n6036), .B (n7642), .Y (y3901) );
  AO21x1_ASAP7_75t_R   g7636( .A1 (n22), .A2 (n17), .B (n3310), .Y (n7644) );
  AO21x1_ASAP7_75t_R   g7637( .A1 (n4129), .A2 (n348), .B (x5), .Y (n7645) );
  OA21x2_ASAP7_75t_R   g7638( .A1 (n7644), .A2 (n7619), .B (n7645), .Y (y3902) );
  AO21x1_ASAP7_75t_R   g7639( .A1 (n466), .A2 (n58), .B (n972), .Y (y3903) );
  NAND2x1_ASAP7_75t_R  g7640( .A (x5), .B (n3310), .Y (n7648) );
  INVx1_ASAP7_75t_R    g7641( .A (n7648), .Y (n7649) );
  AO21x1_ASAP7_75t_R   g7642( .A1 (n15), .A2 (x5), .B (n325), .Y (n7650) );
  INVx1_ASAP7_75t_R    g7643( .A (n7650), .Y (n7651) );
  OR3x1_ASAP7_75t_R    g7644( .A (n7649), .B (n4188), .C (n7651), .Y (y3904) );
  INVx1_ASAP7_75t_R    g7645( .A (n4439), .Y (n7653) );
  NAND2x1_ASAP7_75t_R  g7646( .A (x5), .B (n7653), .Y (n7654) );
  OA33x2_ASAP7_75t_R   g7647( .A1 (n211), .A2 (n421), .A3 (n3637), .B1 (n164), .B2 (n7654), .B3 (n671), .Y (y3905) );
  NAND2x1_ASAP7_75t_R  g7648( .A (n4439), .B (n3001), .Y (n7656) );
  AO21x1_ASAP7_75t_R   g7649( .A1 (n5065), .A2 (n7656), .B (n3568), .Y (y3906) );
  NAND2x1_ASAP7_75t_R  g7650( .A (n388), .B (n72), .Y (n7658) );
  AO32x1_ASAP7_75t_R   g7651( .A1 (n388), .A2 (n72), .A3 (n4439), .B1 (n7653), .B2 (n7658), .Y (y3907) );
  AO21x1_ASAP7_75t_R   g7652( .A1 (y9), .A2 (n856), .B (n143), .Y (n7660) );
  AND2x2_ASAP7_75t_R   g7653( .A (n7660), .B (n2116), .Y (y3908) );
  AO32x1_ASAP7_75t_R   g7654( .A1 (n22), .A2 (n397), .A3 (n5963), .B1 (x4), .B2 (n3193), .Y (y3909) );
  AND3x1_ASAP7_75t_R   g7655( .A (y3198), .B (n3797), .C (n299), .Y (y3910) );
  AND3x1_ASAP7_75t_R   g7656( .A (y3758), .B (n72), .C (n137), .Y (n7664) );
  AO21x1_ASAP7_75t_R   g7657( .A1 (n3493), .A2 (n396), .B (n7664), .Y (n7665) );
  OR3x1_ASAP7_75t_R    g7658( .A (n7665), .B (n3568), .C (n628), .Y (y3911) );
  AO21x1_ASAP7_75t_R   g7659( .A1 (n180), .A2 (n56), .B (y1201), .Y (y3912) );
  AND3x1_ASAP7_75t_R   g7660( .A (n2323), .B (n219), .C (n64), .Y (y3913) );
  OA211x2_ASAP7_75t_R  g7661( .A1 (n7658), .A2 (n7653), .B (n3718), .C (n1265), .Y (n7669) );
  INVx1_ASAP7_75t_R    g7662( .A (n7669), .Y (y3914) );
  NAND2x1_ASAP7_75t_R  g7663( .A (n99), .B (n692), .Y (y3915) );
  AND2x2_ASAP7_75t_R   g7664( .A (n2322), .B (n2338), .Y (y3916) );
  INVx1_ASAP7_75t_R    g7665( .A (n3237), .Y (n7673) );
  AND3x1_ASAP7_75t_R   g7666( .A (n7673), .B (n360), .C (n319), .Y (n7674) );
  INVx1_ASAP7_75t_R    g7667( .A (n7674), .Y (n7675) );
  AND2x2_ASAP7_75t_R   g7668( .A (n7675), .B (n4317), .Y (y3917) );
  AND2x2_ASAP7_75t_R   g7669( .A (n3968), .B (n4108), .Y (y3918) );
  OA21x2_ASAP7_75t_R   g7670( .A1 (n3548), .A2 (n3896), .B (n4089), .Y (y3919) );
  AND3x1_ASAP7_75t_R   g7671( .A (n72), .B (n22), .C (x5), .Y (n7679) );
  OR3x1_ASAP7_75t_R    g7672( .A (n7679), .B (n4915), .C (n628), .Y (y3920) );
  AND3x1_ASAP7_75t_R   g7673( .A (n3469), .B (n3685), .C (x5), .Y (n7681) );
  AO21x1_ASAP7_75t_R   g7674( .A1 (n3183), .A2 (n4924), .B (n7681), .Y (y3921) );
  NOR2x1_ASAP7_75t_R   g7675( .A (x5), .B (n7209), .Y (y3922) );
  AO21x1_ASAP7_75t_R   g7676( .A1 (x2), .A2 (n22), .B (n369), .Y (n7684) );
  AO21x1_ASAP7_75t_R   g7677( .A1 (n7684), .A2 (n3469), .B (n3333), .Y (y3923) );
  OA21x2_ASAP7_75t_R   g7678( .A1 (n3298), .A2 (n5108), .B (n4109), .Y (y3924) );
  AO21x1_ASAP7_75t_R   g7679( .A1 (n17), .A2 (n22), .B (n756), .Y (n7687) );
  AO21x1_ASAP7_75t_R   g7680( .A1 (n7687), .A2 (n7588), .B (n3566), .Y (y3925) );
  OR3x1_ASAP7_75t_R    g7681( .A (n7679), .B (n4915), .C (n3960), .Y (y3926) );
  AO21x1_ASAP7_75t_R   g7682( .A1 (n4755), .A2 (n5090), .B (n164), .Y (y3927) );
  AND2x2_ASAP7_75t_R   g7683( .A (n3987), .B (y1890), .Y (y3928) );
  NOR2x1_ASAP7_75t_R   g7684( .A (n12), .B (n1644), .Y (n7692) );
  OR3x1_ASAP7_75t_R    g7685( .A (n7692), .B (n791), .C (n495), .Y (y3929) );
  INVx1_ASAP7_75t_R    g7686( .A (n6504), .Y (n7694) );
  AO21x1_ASAP7_75t_R   g7687( .A1 (n7694), .A2 (x3), .B (n4981), .Y (y3930) );
  AND2x2_ASAP7_75t_R   g7688( .A (n1283), .B (n1326), .Y (y3931) );
  AO21x1_ASAP7_75t_R   g7689( .A1 (x2), .A2 (n3338), .B (n7658), .Y (y3932) );
  AO21x1_ASAP7_75t_R   g7690( .A1 (n17), .A2 (n310), .B (n300), .Y (n7698) );
  AO21x1_ASAP7_75t_R   g7691( .A1 (n7698), .A2 (n299), .B (n628), .Y (y3933) );
  NOR2x1_ASAP7_75t_R   g7692( .A (n4240), .B (n5251), .Y (y3934) );
  NOR2x1_ASAP7_75t_R   g7693( .A (n918), .B (n6040), .Y (y3935) );
  OA21x2_ASAP7_75t_R   g7694( .A1 (x3), .A2 (n308), .B (n6871), .Y (y3936) );
  AO21x1_ASAP7_75t_R   g7695( .A1 (n1158), .A2 (n97), .B (n3278), .Y (y3937) );
  AO21x1_ASAP7_75t_R   g7696( .A1 (n15), .A2 (y2079), .B (n3027), .Y (n7704) );
  AO21x1_ASAP7_75t_R   g7697( .A1 (n7704), .A2 (n388), .B (n17), .Y (n7705) );
  NAND2x1_ASAP7_75t_R  g7698( .A (n4216), .B (n7705), .Y (y3938) );
  AO21x1_ASAP7_75t_R   g7699( .A1 (n7654), .A2 (n4789), .B (n3333), .Y (y3941) );
  INVx1_ASAP7_75t_R    g7700( .A (n4619), .Y (n7708) );
  AO21x1_ASAP7_75t_R   g7701( .A1 (n7708), .A2 (n15), .B (n5568), .Y (n7709) );
  OR3x1_ASAP7_75t_R    g7702( .A (n392), .B (n15), .C (n17), .Y (n7710) );
  NAND2x1_ASAP7_75t_R  g7703( .A (n7709), .B (n7710), .Y (y3942) );
  AO21x1_ASAP7_75t_R   g7704( .A1 (n3677), .A2 (n3678), .B (y1802), .Y (n7712) );
  INVx1_ASAP7_75t_R    g7705( .A (n7712), .Y (y3943) );
  AO32x1_ASAP7_75t_R   g7706( .A1 (n15), .A2 (n348), .A3 (x5), .B1 (n2980), .B2 (y3808), .Y (y3944) );
  BUFx2_ASAP7_75t_R    g7707( .A (x0), .Y (y3945) );
  NAND2x1_ASAP7_75t_R  g7708( .A (x5), .B (n5243), .Y (n7716) );
  AO21x1_ASAP7_75t_R   g7709( .A1 (n684), .A2 (n7716), .B (n5117), .Y (y3946) );
  NAND2x1_ASAP7_75t_R  g7710( .A (n3148), .B (n430), .Y (n7718) );
  OR3x1_ASAP7_75t_R    g7711( .A (n418), .B (n12), .C (x1), .Y (n7719) );
  OA21x2_ASAP7_75t_R   g7712( .A1 (n7718), .A2 (n606), .B (n7719), .Y (y3947) );
  NOR2x1_ASAP7_75t_R   g7713( .A (n4631), .B (n7107), .Y (y3948) );
  AND3x1_ASAP7_75t_R   g7714( .A (n76), .B (x5), .C (x4), .Y (n7722) );
  INVx1_ASAP7_75t_R    g7715( .A (n7722), .Y (y3949) );
  NOR2x1_ASAP7_75t_R   g7716( .A (n12), .B (n690), .Y (y3950) );
  AND3x1_ASAP7_75t_R   g7717( .A (y863), .B (x3), .C (x2), .Y (y3951) );
  AND3x1_ASAP7_75t_R   g7718( .A (n466), .B (n219), .C (y2079), .Y (y3952) );
  AO21x1_ASAP7_75t_R   g7719( .A1 (y2079), .A2 (n3377), .B (n4420), .Y (y3953) );
  AO21x1_ASAP7_75t_R   g7720( .A1 (n16), .A2 (n12), .B (n76), .Y (n7728) );
  AND2x2_ASAP7_75t_R   g7721( .A (n7728), .B (n2922), .Y (y3954) );
  OR3x1_ASAP7_75t_R    g7722( .A (n529), .B (n1082), .C (n12), .Y (n7730) );
  AND2x2_ASAP7_75t_R   g7723( .A (n7730), .B (n3880), .Y (y3955) );
  AND2x2_ASAP7_75t_R   g7724( .A (n4789), .B (n3919), .Y (y3956) );
  AND3x1_ASAP7_75t_R   g7725( .A (n6068), .B (n137), .C (n63), .Y (y3957) );
  OA21x2_ASAP7_75t_R   g7726( .A1 (n221), .A2 (n76), .B (n2922), .Y (y3958) );
  AO21x1_ASAP7_75t_R   g7727( .A1 (n15), .A2 (n5764), .B (y2916), .Y (y3959) );
  OA21x2_ASAP7_75t_R   g7728( .A1 (n2841), .A2 (n81), .B (x0), .Y (y3960) );
  AO21x1_ASAP7_75t_R   g7729( .A1 (n189), .A2 (y2079), .B (n337), .Y (y3961) );
  OA21x2_ASAP7_75t_R   g7730( .A1 (n81), .A2 (n2841), .B (n219), .Y (y3962) );
  INVx1_ASAP7_75t_R    g7731( .A (n851), .Y (n7739) );
  AO21x1_ASAP7_75t_R   g7732( .A1 (n7739), .A2 (n1373), .B (n143), .Y (y3964) );
  OA21x2_ASAP7_75t_R   g7733( .A1 (n5978), .A2 (x3), .B (n4099), .Y (y3965) );
  NAND2x1_ASAP7_75t_R  g7734( .A (n15), .B (n2256), .Y (n7742) );
  OA211x2_ASAP7_75t_R  g7735( .A1 (n137), .A2 (n227), .B (n7742), .C (n5393), .Y (y3966) );
  AO21x1_ASAP7_75t_R   g7736( .A1 (n4824), .A2 (n419), .B (x0), .Y (y3967) );
  AO21x1_ASAP7_75t_R   g7737( .A1 (n3164), .A2 (n52), .B (x0), .Y (y3969) );
  AO21x1_ASAP7_75t_R   g7738( .A1 (n5030), .A2 (n3284), .B (n3719), .Y (y3970) );
  AO21x1_ASAP7_75t_R   g7739( .A1 (x3), .A2 (n16), .B (n1469), .Y (n7747) );
  INVx1_ASAP7_75t_R    g7740( .A (n7747), .Y (n7748) );
  OA21x2_ASAP7_75t_R   g7741( .A1 (n7748), .A2 (n2889), .B (n152), .Y (y3971) );
  AOI22x1_ASAP7_75t_R  g7742( .A1 (n2583), .A2 (n622), .B1 (x3), .B2 (n1301), .Y (y3972) );
  NAND2x1_ASAP7_75t_R  g7743( .A (n30), .B (y3852), .Y (n7751) );
  NAND2x1_ASAP7_75t_R  g7744( .A (x1), .B (n386), .Y (n7752) );
  AO21x1_ASAP7_75t_R   g7745( .A1 (n7751), .A2 (n7752), .B (n914), .Y (y3973) );
  AND3x1_ASAP7_75t_R   g7746( .A (n2754), .B (n236), .C (n171), .Y (y3974) );
  AO21x1_ASAP7_75t_R   g7747( .A1 (n3850), .A2 (n556), .B (n1277), .Y (y3975) );
  AO21x1_ASAP7_75t_R   g7748( .A1 (n17), .A2 (x2), .B (y863), .Y (n7756) );
  AND3x1_ASAP7_75t_R   g7749( .A (n7756), .B (n228), .C (n72), .Y (n7757) );
  NAND2x1_ASAP7_75t_R  g7750( .A (x1), .B (n70), .Y (n7758) );
  AND2x2_ASAP7_75t_R   g7751( .A (n7757), .B (n7758), .Y (y3976) );
  NAND2x1_ASAP7_75t_R  g7752( .A (n1676), .B (n5210), .Y (y3977) );
  AO21x1_ASAP7_75t_R   g7753( .A1 (n28), .A2 (n352), .B (x3), .Y (n7761) );
  AND2x2_ASAP7_75t_R   g7754( .A (n922), .B (n7761), .Y (y3978) );
  NAND2x1_ASAP7_75t_R  g7755( .A (x0), .B (n151), .Y (n7763) );
  AND3x1_ASAP7_75t_R   g7756( .A (n7763), .B (n3721), .C (n113), .Y (y3979) );
  AND2x2_ASAP7_75t_R   g7757( .A (n3455), .B (x0), .Y (y3981) );
  OA22x2_ASAP7_75t_R   g7758( .A1 (n2583), .A2 (n4602), .B1 (n5790), .B2 (n45), .Y (y3982) );
  AO21x1_ASAP7_75t_R   g7759( .A1 (y9), .A2 (n17), .B (n2169), .Y (n7767) );
  AND2x2_ASAP7_75t_R   g7760( .A (n7763), .B (n7767), .Y (y3983) );
endmodule
